module ShiftRegister(
  input          clock,
  input  [127:0] io_input,
  input          io_enable,
  input          io_rev,
  input          io_cyc,
  input          io_tap,
  output [127:0] io_output_0,
  output [127:0] io_output_1,
  output [127:0] io_output_2,
  output [127:0] io_output_3,
  output [127:0] io_output_4,
  output [127:0] io_output_5,
  output [127:0] io_output_6,
  output [127:0] io_output_7,
  output [127:0] io_output_8,
  output [127:0] io_output_9,
  output [127:0] io_output_10,
  output [127:0] io_output_11,
  output [127:0] io_output_12,
  output [127:0] io_output_13,
  output [127:0] io_output_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] reg_0; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_1; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_2; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_3; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_4; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_5; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_6; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_7; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_8; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_9; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_10; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_11; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_12; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_13; // @[ShiftRegister.scala 34:18]
  reg [127:0] reg_14; // @[ShiftRegister.scala 34:18]
  wire [2:0] _T = io_tap ? 3'h0 : 3'h4; // @[ShiftRegister.scala 42:36]
  wire [3:0] _GEN_75 = {{1'd0}, _T}; // @[ShiftRegister.scala 42:26]
  assign io_output_0 = reg_0; // @[ShiftRegister.scala 53:15]
  assign io_output_1 = reg_1; // @[ShiftRegister.scala 53:15]
  assign io_output_2 = reg_2; // @[ShiftRegister.scala 53:15]
  assign io_output_3 = reg_3; // @[ShiftRegister.scala 53:15]
  assign io_output_4 = reg_4; // @[ShiftRegister.scala 53:15]
  assign io_output_5 = reg_5; // @[ShiftRegister.scala 53:15]
  assign io_output_6 = reg_6; // @[ShiftRegister.scala 53:15]
  assign io_output_7 = reg_7; // @[ShiftRegister.scala 53:15]
  assign io_output_8 = reg_8; // @[ShiftRegister.scala 53:15]
  assign io_output_9 = reg_9; // @[ShiftRegister.scala 53:15]
  assign io_output_10 = reg_10; // @[ShiftRegister.scala 53:15]
  assign io_output_11 = reg_11; // @[ShiftRegister.scala 53:15]
  assign io_output_12 = reg_12; // @[ShiftRegister.scala 53:15]
  assign io_output_13 = reg_13; // @[ShiftRegister.scala 53:15]
  assign io_output_14 = reg_14; // @[ShiftRegister.scala 53:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  reg_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  reg_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  reg_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  reg_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  reg_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  reg_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  reg_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  reg_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  reg_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  reg_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  reg_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  reg_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  reg_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  reg_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  reg_14 = _RAND_14[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_enable) begin
      if (io_rev) begin
        reg_0 <= reg_1;
      end else if (io_cyc) begin
        if (3'h0 == _T) begin
          reg_0 <= reg_14;
        end
      end else begin
        reg_0 <= io_input;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_1 <= reg_2;
      end else if (io_cyc) begin
        if (3'h1 == _T) begin
          reg_1 <= reg_14;
        end else begin
          reg_1 <= reg_0;
        end
      end else begin
        reg_1 <= reg_0;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_2 <= reg_3;
      end else if (io_cyc) begin
        if (3'h2 == _T) begin
          reg_2 <= reg_14;
        end else begin
          reg_2 <= reg_1;
        end
      end else begin
        reg_2 <= reg_1;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_3 <= reg_4;
      end else if (io_cyc) begin
        if (3'h3 == _T) begin
          reg_3 <= reg_14;
        end else begin
          reg_3 <= reg_2;
        end
      end else begin
        reg_3 <= reg_2;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_4 <= reg_5;
      end else if (io_cyc) begin
        if (3'h4 == _T) begin
          reg_4 <= reg_14;
        end else begin
          reg_4 <= reg_3;
        end
      end else begin
        reg_4 <= reg_3;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_5 <= reg_6;
      end else if (io_cyc) begin
        if (3'h5 == _T) begin
          reg_5 <= reg_14;
        end else begin
          reg_5 <= reg_4;
        end
      end else begin
        reg_5 <= reg_4;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_6 <= reg_7;
      end else if (io_cyc) begin
        if (3'h6 == _T) begin
          reg_6 <= reg_14;
        end else begin
          reg_6 <= reg_5;
        end
      end else begin
        reg_6 <= reg_5;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_7 <= reg_8;
      end else if (io_cyc) begin
        if (3'h7 == _T) begin
          reg_7 <= reg_14;
        end else begin
          reg_7 <= reg_6;
        end
      end else begin
        reg_7 <= reg_6;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_8 <= reg_9;
      end else if (io_cyc) begin
        if (4'h8 == _GEN_75) begin
          reg_8 <= reg_14;
        end else begin
          reg_8 <= reg_7;
        end
      end else begin
        reg_8 <= reg_7;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_9 <= reg_10;
      end else if (io_cyc) begin
        if (4'h9 == _GEN_75) begin
          reg_9 <= reg_14;
        end else begin
          reg_9 <= reg_8;
        end
      end else begin
        reg_9 <= reg_8;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_10 <= reg_11;
      end else if (io_cyc) begin
        if (4'ha == _GEN_75) begin
          reg_10 <= reg_14;
        end else begin
          reg_10 <= reg_9;
        end
      end else begin
        reg_10 <= reg_9;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_11 <= reg_12;
      end else if (io_cyc) begin
        if (4'hb == _GEN_75) begin
          reg_11 <= reg_14;
        end else begin
          reg_11 <= reg_10;
        end
      end else begin
        reg_11 <= reg_10;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_12 <= reg_13;
      end else if (io_cyc) begin
        if (4'hc == _GEN_75) begin
          reg_12 <= reg_14;
        end else begin
          reg_12 <= reg_11;
        end
      end else begin
        reg_12 <= reg_11;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        reg_13 <= reg_14;
      end else if (io_cyc) begin
        if (4'hd == _GEN_75) begin
          reg_13 <= reg_14;
        end else begin
          reg_13 <= reg_12;
        end
      end else begin
        reg_13 <= reg_12;
      end
    end
    if (io_enable) begin
      if (io_rev) begin
        if (!(4'he == _GEN_75)) begin
          if (4'hd == _GEN_75) begin
            reg_14 <= reg_13;
          end else if (4'hc == _GEN_75) begin
            reg_14 <= reg_12;
          end else if (4'hb == _GEN_75) begin
            reg_14 <= reg_11;
          end else if (4'ha == _GEN_75) begin
            reg_14 <= reg_10;
          end else if (4'h9 == _GEN_75) begin
            reg_14 <= reg_9;
          end else if (4'h8 == _GEN_75) begin
            reg_14 <= reg_8;
          end else if (3'h7 == _T) begin
            reg_14 <= reg_7;
          end else if (3'h6 == _T) begin
            reg_14 <= reg_6;
          end else if (3'h5 == _T) begin
            reg_14 <= reg_5;
          end else if (3'h4 == _T) begin
            reg_14 <= reg_4;
          end else if (3'h3 == _T) begin
            reg_14 <= reg_3;
          end else if (3'h2 == _T) begin
            reg_14 <= reg_2;
          end else if (3'h1 == _T) begin
            reg_14 <= reg_1;
          end else begin
            reg_14 <= reg_0;
          end
        end
      end else if (io_cyc) begin
        if (!(4'he == _GEN_75)) begin
          reg_14 <= reg_13;
        end
      end else begin
        reg_14 <= reg_13;
      end
    end
  end
endmodule
module MixColsModule(
  input  [7:0] io_in_0_0,
  input  [7:0] io_in_0_1,
  input  [7:0] io_in_0_2,
  input  [7:0] io_in_0_3,
  input  [7:0] io_in_1_0,
  input  [7:0] io_in_1_1,
  input  [7:0] io_in_1_2,
  input  [7:0] io_in_1_3,
  input  [7:0] io_in_2_0,
  input  [7:0] io_in_2_1,
  input  [7:0] io_in_2_2,
  input  [7:0] io_in_2_3,
  input  [7:0] io_in_3_0,
  input  [7:0] io_in_3_1,
  input  [7:0] io_in_3_2,
  input  [7:0] io_in_3_3,
  output [7:0] io_out_0_0,
  output [7:0] io_out_0_1,
  output [7:0] io_out_0_2,
  output [7:0] io_out_0_3,
  output [7:0] io_out_1_0,
  output [7:0] io_out_1_1,
  output [7:0] io_out_1_2,
  output [7:0] io_out_1_3,
  output [7:0] io_out_2_0,
  output [7:0] io_out_2_1,
  output [7:0] io_out_2_2,
  output [7:0] io_out_2_3,
  output [7:0] io_out_3_0,
  output [7:0] io_out_3_1,
  output [7:0] io_out_3_2,
  output [7:0] io_out_3_3
);
  wire [7:0] _T = io_in_0_0 ^ io_in_0_1; // @[AesComponents.scala 30:29]
  wire [7:0] _T_1 = _T ^ io_in_0_2; // @[AesComponents.scala 30:43]
  wire [7:0] _T_2 = _T_1 ^ io_in_0_3; // @[AesComponents.scala 30:57]
  wire [7:0] _T_3 = io_in_0_0 ^ _T_2; // @[AesComponents.scala 31:37]
  wire [7:0] _T_5 = _T & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_6 = _T_5 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_7 = {_T, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_8 = _T_7 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_9 = _T_8 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_11 = _T_6 ? _T_9 : _T_7; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_0 = {{1'd0}, _T_3}; // @[AesComponents.scala 31:41]
  wire [8:0] _T_12 = _GEN_0 ^ _T_11; // @[AesComponents.scala 31:41]
  wire [7:0] _T_13 = io_in_0_1 ^ _T_2; // @[AesComponents.scala 32:37]
  wire [7:0] _T_14 = io_in_0_1 ^ io_in_0_2; // @[AesComponents.scala 32:64]
  wire [7:0] _T_15 = _T_14 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_16 = _T_15 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_17 = {_T_14, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_18 = _T_17 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_19 = _T_18 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_21 = _T_16 ? _T_19 : _T_17; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_1 = {{1'd0}, _T_13}; // @[AesComponents.scala 32:41]
  wire [8:0] _T_22 = _GEN_1 ^ _T_21; // @[AesComponents.scala 32:41]
  wire [7:0] _T_23 = io_in_0_2 ^ _T_2; // @[AesComponents.scala 33:37]
  wire [7:0] _T_24 = io_in_0_2 ^ io_in_0_3; // @[AesComponents.scala 33:64]
  wire [7:0] _T_25 = _T_24 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_26 = _T_25 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_27 = {_T_24, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_28 = _T_27 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_29 = _T_28 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_31 = _T_26 ? _T_29 : _T_27; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_2 = {{1'd0}, _T_23}; // @[AesComponents.scala 33:41]
  wire [8:0] _T_32 = _GEN_2 ^ _T_31; // @[AesComponents.scala 33:41]
  wire [7:0] _T_33 = io_in_0_3 ^ _T_2; // @[AesComponents.scala 34:37]
  wire [7:0] _T_34 = io_in_0_3 ^ io_in_0_0; // @[AesComponents.scala 34:64]
  wire [7:0] _T_35 = _T_34 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_36 = _T_35 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_37 = {_T_34, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_38 = _T_37 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_39 = _T_38 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_41 = _T_36 ? _T_39 : _T_37; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_3 = {{1'd0}, _T_33}; // @[AesComponents.scala 34:41]
  wire [8:0] _T_42 = _GEN_3 ^ _T_41; // @[AesComponents.scala 34:41]
  wire [7:0] _T_43 = io_in_1_0 ^ io_in_1_1; // @[AesComponents.scala 30:29]
  wire [7:0] _T_44 = _T_43 ^ io_in_1_2; // @[AesComponents.scala 30:43]
  wire [7:0] _T_45 = _T_44 ^ io_in_1_3; // @[AesComponents.scala 30:57]
  wire [7:0] _T_46 = io_in_1_0 ^ _T_45; // @[AesComponents.scala 31:37]
  wire [7:0] _T_48 = _T_43 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_49 = _T_48 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_50 = {_T_43, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_51 = _T_50 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_52 = _T_51 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_54 = _T_49 ? _T_52 : _T_50; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_4 = {{1'd0}, _T_46}; // @[AesComponents.scala 31:41]
  wire [8:0] _T_55 = _GEN_4 ^ _T_54; // @[AesComponents.scala 31:41]
  wire [7:0] _T_56 = io_in_1_1 ^ _T_45; // @[AesComponents.scala 32:37]
  wire [7:0] _T_57 = io_in_1_1 ^ io_in_1_2; // @[AesComponents.scala 32:64]
  wire [7:0] _T_58 = _T_57 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_59 = _T_58 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_60 = {_T_57, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_61 = _T_60 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_62 = _T_61 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_64 = _T_59 ? _T_62 : _T_60; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_5 = {{1'd0}, _T_56}; // @[AesComponents.scala 32:41]
  wire [8:0] _T_65 = _GEN_5 ^ _T_64; // @[AesComponents.scala 32:41]
  wire [7:0] _T_66 = io_in_1_2 ^ _T_45; // @[AesComponents.scala 33:37]
  wire [7:0] _T_67 = io_in_1_2 ^ io_in_1_3; // @[AesComponents.scala 33:64]
  wire [7:0] _T_68 = _T_67 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_69 = _T_68 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_70 = {_T_67, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_71 = _T_70 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_72 = _T_71 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_74 = _T_69 ? _T_72 : _T_70; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_6 = {{1'd0}, _T_66}; // @[AesComponents.scala 33:41]
  wire [8:0] _T_75 = _GEN_6 ^ _T_74; // @[AesComponents.scala 33:41]
  wire [7:0] _T_76 = io_in_1_3 ^ _T_45; // @[AesComponents.scala 34:37]
  wire [7:0] _T_77 = io_in_1_3 ^ io_in_1_0; // @[AesComponents.scala 34:64]
  wire [7:0] _T_78 = _T_77 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_79 = _T_78 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_80 = {_T_77, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_81 = _T_80 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_82 = _T_81 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_84 = _T_79 ? _T_82 : _T_80; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_7 = {{1'd0}, _T_76}; // @[AesComponents.scala 34:41]
  wire [8:0] _T_85 = _GEN_7 ^ _T_84; // @[AesComponents.scala 34:41]
  wire [7:0] _T_86 = io_in_2_0 ^ io_in_2_1; // @[AesComponents.scala 30:29]
  wire [7:0] _T_87 = _T_86 ^ io_in_2_2; // @[AesComponents.scala 30:43]
  wire [7:0] _T_88 = _T_87 ^ io_in_2_3; // @[AesComponents.scala 30:57]
  wire [7:0] _T_89 = io_in_2_0 ^ _T_88; // @[AesComponents.scala 31:37]
  wire [7:0] _T_91 = _T_86 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_92 = _T_91 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_93 = {_T_86, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_94 = _T_93 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_95 = _T_94 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_97 = _T_92 ? _T_95 : _T_93; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_8 = {{1'd0}, _T_89}; // @[AesComponents.scala 31:41]
  wire [8:0] _T_98 = _GEN_8 ^ _T_97; // @[AesComponents.scala 31:41]
  wire [7:0] _T_99 = io_in_2_1 ^ _T_88; // @[AesComponents.scala 32:37]
  wire [7:0] _T_100 = io_in_2_1 ^ io_in_2_2; // @[AesComponents.scala 32:64]
  wire [7:0] _T_101 = _T_100 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_102 = _T_101 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_103 = {_T_100, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_104 = _T_103 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_105 = _T_104 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_107 = _T_102 ? _T_105 : _T_103; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_9 = {{1'd0}, _T_99}; // @[AesComponents.scala 32:41]
  wire [8:0] _T_108 = _GEN_9 ^ _T_107; // @[AesComponents.scala 32:41]
  wire [7:0] _T_109 = io_in_2_2 ^ _T_88; // @[AesComponents.scala 33:37]
  wire [7:0] _T_110 = io_in_2_2 ^ io_in_2_3; // @[AesComponents.scala 33:64]
  wire [7:0] _T_111 = _T_110 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_112 = _T_111 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_113 = {_T_110, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_114 = _T_113 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_115 = _T_114 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_117 = _T_112 ? _T_115 : _T_113; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_10 = {{1'd0}, _T_109}; // @[AesComponents.scala 33:41]
  wire [8:0] _T_118 = _GEN_10 ^ _T_117; // @[AesComponents.scala 33:41]
  wire [7:0] _T_119 = io_in_2_3 ^ _T_88; // @[AesComponents.scala 34:37]
  wire [7:0] _T_120 = io_in_2_3 ^ io_in_2_0; // @[AesComponents.scala 34:64]
  wire [7:0] _T_121 = _T_120 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_122 = _T_121 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_123 = {_T_120, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_124 = _T_123 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_125 = _T_124 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_127 = _T_122 ? _T_125 : _T_123; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_11 = {{1'd0}, _T_119}; // @[AesComponents.scala 34:41]
  wire [8:0] _T_128 = _GEN_11 ^ _T_127; // @[AesComponents.scala 34:41]
  wire [7:0] _T_129 = io_in_3_0 ^ io_in_3_1; // @[AesComponents.scala 30:29]
  wire [7:0] _T_130 = _T_129 ^ io_in_3_2; // @[AesComponents.scala 30:43]
  wire [7:0] _T_131 = _T_130 ^ io_in_3_3; // @[AesComponents.scala 30:57]
  wire [7:0] _T_132 = io_in_3_0 ^ _T_131; // @[AesComponents.scala 31:37]
  wire [7:0] _T_134 = _T_129 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_135 = _T_134 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_136 = {_T_129, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_137 = _T_136 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_138 = _T_137 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_140 = _T_135 ? _T_138 : _T_136; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_12 = {{1'd0}, _T_132}; // @[AesComponents.scala 31:41]
  wire [8:0] _T_141 = _GEN_12 ^ _T_140; // @[AesComponents.scala 31:41]
  wire [7:0] _T_142 = io_in_3_1 ^ _T_131; // @[AesComponents.scala 32:37]
  wire [7:0] _T_143 = io_in_3_1 ^ io_in_3_2; // @[AesComponents.scala 32:64]
  wire [7:0] _T_144 = _T_143 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_145 = _T_144 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_146 = {_T_143, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_147 = _T_146 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_148 = _T_147 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_150 = _T_145 ? _T_148 : _T_146; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_13 = {{1'd0}, _T_142}; // @[AesComponents.scala 32:41]
  wire [8:0] _T_151 = _GEN_13 ^ _T_150; // @[AesComponents.scala 32:41]
  wire [7:0] _T_152 = io_in_3_2 ^ _T_131; // @[AesComponents.scala 33:37]
  wire [7:0] _T_153 = io_in_3_2 ^ io_in_3_3; // @[AesComponents.scala 33:64]
  wire [7:0] _T_154 = _T_153 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_155 = _T_154 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_156 = {_T_153, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_157 = _T_156 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_158 = _T_157 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_160 = _T_155 ? _T_158 : _T_156; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_14 = {{1'd0}, _T_152}; // @[AesComponents.scala 33:41]
  wire [8:0] _T_161 = _GEN_14 ^ _T_160; // @[AesComponents.scala 33:41]
  wire [7:0] _T_162 = io_in_3_3 ^ _T_131; // @[AesComponents.scala 34:37]
  wire [7:0] _T_163 = io_in_3_3 ^ io_in_3_0; // @[AesComponents.scala 34:64]
  wire [7:0] _T_164 = _T_163 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_165 = _T_164 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_166 = {_T_163, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_167 = _T_166 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_168 = _T_167 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_170 = _T_165 ? _T_168 : _T_166; // @[AesComponents.scala 88:38]
  wire [8:0] _GEN_15 = {{1'd0}, _T_162}; // @[AesComponents.scala 34:41]
  wire [8:0] _T_171 = _GEN_15 ^ _T_170; // @[AesComponents.scala 34:41]
  assign io_out_0_0 = _T_12[7:0]; // @[AesComponents.scala 31:22]
  assign io_out_0_1 = _T_22[7:0]; // @[AesComponents.scala 32:22]
  assign io_out_0_2 = _T_32[7:0]; // @[AesComponents.scala 33:22]
  assign io_out_0_3 = _T_42[7:0]; // @[AesComponents.scala 34:22]
  assign io_out_1_0 = _T_55[7:0]; // @[AesComponents.scala 31:22]
  assign io_out_1_1 = _T_65[7:0]; // @[AesComponents.scala 32:22]
  assign io_out_1_2 = _T_75[7:0]; // @[AesComponents.scala 33:22]
  assign io_out_1_3 = _T_85[7:0]; // @[AesComponents.scala 34:22]
  assign io_out_2_0 = _T_98[7:0]; // @[AesComponents.scala 31:22]
  assign io_out_2_1 = _T_108[7:0]; // @[AesComponents.scala 32:22]
  assign io_out_2_2 = _T_118[7:0]; // @[AesComponents.scala 33:22]
  assign io_out_2_3 = _T_128[7:0]; // @[AesComponents.scala 34:22]
  assign io_out_3_0 = _T_141[7:0]; // @[AesComponents.scala 31:22]
  assign io_out_3_1 = _T_151[7:0]; // @[AesComponents.scala 32:22]
  assign io_out_3_2 = _T_161[7:0]; // @[AesComponents.scala 33:22]
  assign io_out_3_3 = _T_171[7:0]; // @[AesComponents.scala 34:22]
endmodule
module AesEncrypt(
  input          clock,
  input          reset,
  input  [127:0] io_dataIn,
  input  [127:0] io_ivIn,
  input          io_dataValid,
  input  [7:0]   io_keys_0_0_0,
  input  [7:0]   io_keys_0_0_1,
  input  [7:0]   io_keys_0_0_2,
  input  [7:0]   io_keys_0_0_3,
  input  [7:0]   io_keys_0_1_0,
  input  [7:0]   io_keys_0_1_1,
  input  [7:0]   io_keys_0_1_2,
  input  [7:0]   io_keys_0_1_3,
  input  [7:0]   io_keys_0_2_0,
  input  [7:0]   io_keys_0_2_1,
  input  [7:0]   io_keys_0_2_2,
  input  [7:0]   io_keys_0_2_3,
  input  [7:0]   io_keys_0_3_0,
  input  [7:0]   io_keys_0_3_1,
  input  [7:0]   io_keys_0_3_2,
  input  [7:0]   io_keys_0_3_3,
  input          io_aes256,
  output         io_shiftCyc,
  output         io_shift,
  output         io_ready,
  output [127:0] io_dataOut,
  output [127:0] io_ivOut,
  output         io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] MixColsModule_io_in_0_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_0_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_0_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_0_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_3; // @[AesComponents.scala 91:35]
  reg [5:0] state; // @[AesEncrypt.scala 54:24]
  wire  _T = state == 6'h0; // @[AesEncrypt.scala 56:24]
  wire  _T_1 = state == 6'h1; // @[AesEncrypt.scala 56:43]
  wire  _T_2 = _T | _T_1; // @[AesEncrypt.scala 56:33]
  wire  _T_3 = state == 6'h1e; // @[AesEncrypt.scala 56:62]
  wire  _T_6 = ~io_ready; // @[AesEncrypt.scala 59:31]
  reg [7:0] matrix_0_0; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_0_1; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_0_2; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_0_3; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_1_0; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_1_1; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_1_2; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_1_3; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_2_0; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_2_1; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_2_2; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_2_3; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_3_0; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_3_1; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_3_2; // @[AesEncrypt.scala 63:21]
  reg [7:0] matrix_3_3; // @[AesEncrypt.scala 63:21]
  wire [63:0] _T_16 = {matrix_2_0,matrix_2_1,matrix_2_2,matrix_2_3,matrix_3_0,matrix_3_1,matrix_3_2,matrix_3_3}; // @[Cat.scala 29:58]
  wire [63:0] _T_23 = {matrix_0_0,matrix_0_1,matrix_0_2,matrix_0_3,matrix_1_0,matrix_1_1,matrix_1_2,matrix_1_3}; // @[Cat.scala 29:58]
  wire [127:0] _T_25 = io_dataIn ^ io_ivIn; // @[AesEncrypt.scala 69:38]
  wire [63:0] _T_32 = {io_keys_0_2_0,io_keys_0_2_1,io_keys_0_2_2,io_keys_0_2_3,io_keys_0_3_0,io_keys_0_3_1,io_keys_0_3_2,io_keys_0_3_3}; // @[Cat.scala 29:58]
  wire [127:0] _T_40 = {io_keys_0_0_0,io_keys_0_0_1,io_keys_0_0_2,io_keys_0_0_3,io_keys_0_1_0,io_keys_0_1_1,io_keys_0_1_2,io_keys_0_1_3,_T_32}; // @[Cat.scala 29:58]
  wire [127:0] _T_41 = _T_25 ^ _T_40; // @[AesEncrypt.scala 69:48]
  wire [7:0] initOut_0_0 = _T_41[127:120]; // @[AesComponents.scala 43:25]
  wire [7:0] initOut_0_1 = _T_41[119:112]; // @[AesComponents.scala 43:45]
  wire [7:0] initOut_0_2 = _T_41[111:104]; // @[AesComponents.scala 43:65]
  wire [7:0] initOut_0_3 = _T_41[103:96]; // @[AesComponents.scala 43:85]
  wire [7:0] initOut_1_0 = _T_41[95:88]; // @[AesComponents.scala 44:25]
  wire [7:0] initOut_1_1 = _T_41[87:80]; // @[AesComponents.scala 44:45]
  wire [7:0] initOut_1_2 = _T_41[79:72]; // @[AesComponents.scala 44:65]
  wire [7:0] initOut_1_3 = _T_41[71:64]; // @[AesComponents.scala 44:85]
  wire [7:0] initOut_2_0 = _T_41[63:56]; // @[AesComponents.scala 45:25]
  wire [7:0] initOut_2_1 = _T_41[55:48]; // @[AesComponents.scala 45:45]
  wire [7:0] initOut_2_2 = _T_41[47:40]; // @[AesComponents.scala 45:65]
  wire [7:0] initOut_2_3 = _T_41[39:32]; // @[AesComponents.scala 45:85]
  wire [7:0] initOut_3_0 = _T_41[31:24]; // @[AesComponents.scala 46:25]
  wire [7:0] initOut_3_1 = _T_41[23:16]; // @[AesComponents.scala 46:45]
  wire [7:0] initOut_3_2 = _T_41[15:8]; // @[AesComponents.scala 46:65]
  wire [7:0] initOut_3_3 = _T_41[7:0]; // @[AesComponents.scala 46:85]
  wire  _T_79 = matrix_0_0[1] ^ matrix_0_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_81 = matrix_0_0[4] ^ matrix_0_0[7]; // @[AesSbox.scala 40:63]
  wire  _T_83 = matrix_0_0[6] ^ matrix_0_0[5]; // @[AesSbox.scala 40:63]
  wire  _T_85 = matrix_0_0[0] ^ _T_83; // @[AesSbox.scala 40:63]
  wire  _T_87 = _T_79 ^ _T_81; // @[AesSbox.scala 40:63]
  wire  _T_89 = matrix_0_0[6] ^ matrix_0_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_91 = matrix_0_0[7] ^ matrix_0_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_93 = _T_79 ^ _T_89; // @[AesSbox.scala 40:63]
  wire  _T_95 = matrix_0_0[1] ^ _T_85; // @[AesSbox.scala 40:63]
  wire  _T_97 = matrix_0_0[4] ^ _T_85; // @[AesSbox.scala 40:63]
  wire  _T_99 = matrix_0_0[0] ^ _T_87; // @[AesSbox.scala 40:63]
  wire  _T_101 = _T_87 ^ _T_89; // @[AesSbox.scala 40:63]
  wire  _T_103 = matrix_0_0[5] ^ matrix_0_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_105 = _T_83 ^ _T_87; // @[AesSbox.scala 40:63]
  wire  _T_107 = matrix_0_0[2] ^ _T_91; // @[AesSbox.scala 40:63]
  wire  _T_109 = matrix_0_0[7] ^ matrix_0_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_111 = matrix_0_0[0] ^ _T_93; // @[AesSbox.scala 40:63]
  wire  _T_113 = matrix_0_0[1] ^ matrix_0_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_115 = _T_81 ^ _T_113; // @[AesSbox.scala 40:63]
  wire  _T_117 = _T_85 ^ _T_107; // @[AesSbox.scala 40:63]
  wire  _T_119 = _T_79 ^ _T_103; // @[AesSbox.scala 40:63]
  wire  _T_121 = matrix_0_0[7] ^ _T_85; // @[AesSbox.scala 40:63]
  wire  _T_123 = _T_119 ^ _T_87; // @[AesSbox.scala 40:63]
  wire  _T_125 = _T_119 ^ _T_91; // @[AesSbox.scala 40:63]
  wire  _T_127 = _T_91 ^ _T_115; // @[AesSbox.scala 40:63]
  wire  _T_129 = _T_109 ^ _T_105; // @[AesSbox.scala 40:63]
  wire  _T_131 = _T_121 ^ _T_111; // @[AesSbox.scala 40:63]
  wire  _T_133 = _T_115 & _T_87; // @[AesSbox.scala 41:63]
  wire  _T_135 = _T_117 & _T_99; // @[AesSbox.scala 41:63]
  wire  _T_137 = _T_101 ^ _T_133; // @[AesSbox.scala 40:63]
  wire  _T_139 = _T_97 & matrix_0_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_141 = _T_139 ^ _T_133; // @[AesSbox.scala 40:63]
  wire  _T_143 = _T_91 & _T_119; // @[AesSbox.scala 41:63]
  wire  _T_145 = _T_95 & _T_85; // @[AesSbox.scala 41:63]
  wire  _T_147 = _T_125 ^ _T_143; // @[AesSbox.scala 40:63]
  wire  _T_149 = _T_121 & _T_111; // @[AesSbox.scala 41:63]
  wire  _T_151 = _T_149 ^ _T_143; // @[AesSbox.scala 40:63]
  wire  _T_153 = _T_81 & _T_93; // @[AesSbox.scala 41:63]
  wire  _T_155 = _T_127 & _T_123; // @[AesSbox.scala 41:63]
  wire  _T_157 = _T_155 ^ _T_153; // @[AesSbox.scala 40:63]
  wire  _T_159 = _T_109 & _T_105; // @[AesSbox.scala 41:63]
  wire  _T_161 = _T_159 ^ _T_153; // @[AesSbox.scala 40:63]
  wire  _T_163 = _T_137 ^ _T_135; // @[AesSbox.scala 40:63]
  wire  _T_165 = _T_141 ^ _T_129; // @[AesSbox.scala 40:63]
  wire  _T_167 = _T_147 ^ _T_145; // @[AesSbox.scala 40:63]
  wire  _T_169 = _T_151 ^ _T_161; // @[AesSbox.scala 40:63]
  wire  _T_171 = _T_163 ^ _T_157; // @[AesSbox.scala 40:63]
  wire  _T_173 = _T_165 ^ _T_161; // @[AesSbox.scala 40:63]
  wire  _T_175 = _T_167 ^ _T_157; // @[AesSbox.scala 40:63]
  wire  _T_177 = _T_169 ^ _T_131; // @[AesSbox.scala 40:63]
  wire  _T_179 = _T_175 ^ _T_177; // @[AesSbox.scala 40:63]
  wire  _T_181 = _T_175 & _T_171; // @[AesSbox.scala 41:63]
  wire  _T_183 = _T_173 ^ _T_181; // @[AesSbox.scala 40:63]
  wire  _T_185 = _T_171 ^ _T_173; // @[AesSbox.scala 40:63]
  wire  _T_187 = _T_177 ^ _T_181; // @[AesSbox.scala 40:63]
  wire  _T_189 = _T_187 & _T_185; // @[AesSbox.scala 41:63]
  wire  _T_191 = _T_183 & _T_179; // @[AesSbox.scala 41:63]
  wire  _T_193 = _T_171 & _T_177; // @[AesSbox.scala 41:63]
  wire  _T_195 = _T_185 & _T_193; // @[AesSbox.scala 41:63]
  wire  _T_197 = _T_185 ^ _T_181; // @[AesSbox.scala 40:63]
  wire  _T_199 = _T_173 & _T_175; // @[AesSbox.scala 41:63]
  wire  _T_201 = _T_179 & _T_199; // @[AesSbox.scala 41:63]
  wire  _T_203 = _T_179 ^ _T_181; // @[AesSbox.scala 40:63]
  wire  _T_205 = _T_173 ^ _T_189; // @[AesSbox.scala 40:63]
  wire  _T_207 = _T_195 ^ _T_197; // @[AesSbox.scala 40:63]
  wire  _T_209 = _T_177 ^ _T_191; // @[AesSbox.scala 40:63]
  wire  _T_211 = _T_201 ^ _T_203; // @[AesSbox.scala 40:63]
  wire  _T_213 = _T_207 ^ _T_211; // @[AesSbox.scala 40:63]
  wire  _T_215 = _T_205 ^ _T_209; // @[AesSbox.scala 40:63]
  wire  _T_217 = _T_205 ^ _T_207; // @[AesSbox.scala 40:63]
  wire  _T_219 = _T_209 ^ _T_211; // @[AesSbox.scala 40:63]
  wire  _T_221 = _T_215 ^ _T_213; // @[AesSbox.scala 40:63]
  wire  _T_223 = _T_219 & _T_87; // @[AesSbox.scala 41:63]
  wire  _T_225 = _T_211 & _T_99; // @[AesSbox.scala 41:63]
  wire  _T_227 = _T_209 & matrix_0_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_229 = _T_217 & _T_119; // @[AesSbox.scala 41:63]
  wire  _T_231 = _T_207 & _T_85; // @[AesSbox.scala 41:63]
  wire  _T_233 = _T_205 & _T_111; // @[AesSbox.scala 41:63]
  wire  _T_235 = _T_215 & _T_93; // @[AesSbox.scala 41:63]
  wire  _T_237 = _T_221 & _T_123; // @[AesSbox.scala 41:63]
  wire  _T_239 = _T_213 & _T_105; // @[AesSbox.scala 41:63]
  wire  _T_241 = _T_219 & _T_115; // @[AesSbox.scala 41:63]
  wire  _T_243 = _T_211 & _T_117; // @[AesSbox.scala 41:63]
  wire  _T_245 = _T_209 & _T_97; // @[AesSbox.scala 41:63]
  wire  _T_247 = _T_217 & _T_91; // @[AesSbox.scala 41:63]
  wire  _T_249 = _T_207 & _T_95; // @[AesSbox.scala 41:63]
  wire  _T_251 = _T_205 & _T_121; // @[AesSbox.scala 41:63]
  wire  _T_253 = _T_215 & _T_81; // @[AesSbox.scala 41:63]
  wire  _T_255 = _T_221 & _T_127; // @[AesSbox.scala 41:63]
  wire  _T_257 = _T_213 & _T_109; // @[AesSbox.scala 41:63]
  wire  _T_259 = _T_253 ^ _T_255; // @[AesSbox.scala 40:63]
  wire  _T_261 = _T_231 ^ _T_243; // @[AesSbox.scala 40:63]
  wire  _T_263 = _T_237 ^ _T_259; // @[AesSbox.scala 40:63]
  wire  _T_265 = _T_241 ^ _T_261; // @[AesSbox.scala 40:63]
  wire  _T_267 = _T_227 ^ _T_247; // @[AesSbox.scala 40:63]
  wire  _T_269 = _T_223 ^ _T_229; // @[AesSbox.scala 40:63]
  wire  _T_271 = _T_259 ^ _T_269; // @[AesSbox.scala 40:63]
  wire  _T_273 = _T_225 ^ _T_265; // @[AesSbox.scala 40:63]
  wire  _T_275 = _T_223 ^ _T_235; // @[AesSbox.scala 40:63]
  wire  _T_277 = _T_233 ^ _T_249; // @[AesSbox.scala 40:63]
  wire  _T_279 = _T_239 ^ _T_251; // @[AesSbox.scala 40:63]
  wire  _T_281 = _T_227 ^ _T_273; // @[AesSbox.scala 40:63]
  wire  _T_283 = _T_267 ^ _T_279; // @[AesSbox.scala 40:63]
  wire  _T_285 = _T_245 ^ _T_261; // @[AesSbox.scala 40:63]
  wire  _T_287 = _T_229 ^ _T_235; // @[AesSbox.scala 40:63]
  wire  _T_289 = _T_265 ^ _T_287; // @[AesSbox.scala 40:63]
  wire  _T_291 = _T_257 ^ _T_283; // @[AesSbox.scala 40:63]
  wire  _T_293 = _T_253 ^ _T_275; // @[AesSbox.scala 40:63]
  wire  _T_295 = _T_267 ^ _T_277; // @[AesSbox.scala 40:63]
  wire  _T_296 = _T_263 ^ _T_289; // @[AesSbox.scala 40:63]
  wire  _T_297 = _T_291 ^ _T_293; // @[AesSbox.scala 42:65]
  wire  _T_298 = ~_T_297; // @[AesSbox.scala 42:51]
  wire  _T_300 = _T_233 ^ _T_259; // @[AesSbox.scala 40:63]
  wire  _T_301 = _T_271 ^ _T_273; // @[AesSbox.scala 40:63]
  wire  _T_302 = _T_281 ^ _T_300; // @[AesSbox.scala 40:63]
  wire  _T_304 = _T_231 ^ _T_247; // @[AesSbox.scala 40:63]
  wire  _T_306 = _T_269 ^ _T_285; // @[AesSbox.scala 40:63]
  wire  _T_307 = _T_271 ^ _T_295; // @[AesSbox.scala 42:65]
  wire  _T_308 = ~_T_307; // @[AesSbox.scala 42:51]
  wire  _T_310 = _T_239 ^ _T_277; // @[AesSbox.scala 40:63]
  wire  _T_312 = _T_304 ^ _T_310; // @[AesSbox.scala 40:63]
  wire  _T_314 = _T_231 ^ _T_275; // @[AesSbox.scala 40:63]
  wire  _T_315 = _T_263 ^ _T_312; // @[AesSbox.scala 42:65]
  wire  _T_316 = ~_T_315; // @[AesSbox.scala 42:51]
  wire  _T_318 = _T_283 ^ _T_306; // @[AesSbox.scala 40:63]
  wire  _T_319 = _T_263 ^ _T_318; // @[AesSbox.scala 40:63]
  wire  _T_321 = _T_273 ^ _T_314; // @[AesSbox.scala 40:63]
  wire  _T_322 = _T_263 ^ _T_321; // @[AesSbox.scala 42:65]
  wire  _T_323 = ~_T_322; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_0_0 = {_T_296,_T_323,_T_298,_T_301,_T_302,_T_319,_T_316,_T_308}; // @[Cat.scala 29:58]
  wire  _T_348 = matrix_0_1[1] ^ matrix_0_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_350 = matrix_0_1[4] ^ matrix_0_1[7]; // @[AesSbox.scala 40:63]
  wire  _T_352 = matrix_0_1[6] ^ matrix_0_1[5]; // @[AesSbox.scala 40:63]
  wire  _T_354 = matrix_0_1[0] ^ _T_352; // @[AesSbox.scala 40:63]
  wire  _T_356 = _T_348 ^ _T_350; // @[AesSbox.scala 40:63]
  wire  _T_358 = matrix_0_1[6] ^ matrix_0_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_360 = matrix_0_1[7] ^ matrix_0_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_362 = _T_348 ^ _T_358; // @[AesSbox.scala 40:63]
  wire  _T_364 = matrix_0_1[1] ^ _T_354; // @[AesSbox.scala 40:63]
  wire  _T_366 = matrix_0_1[4] ^ _T_354; // @[AesSbox.scala 40:63]
  wire  _T_368 = matrix_0_1[0] ^ _T_356; // @[AesSbox.scala 40:63]
  wire  _T_370 = _T_356 ^ _T_358; // @[AesSbox.scala 40:63]
  wire  _T_372 = matrix_0_1[5] ^ matrix_0_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_374 = _T_352 ^ _T_356; // @[AesSbox.scala 40:63]
  wire  _T_376 = matrix_0_1[2] ^ _T_360; // @[AesSbox.scala 40:63]
  wire  _T_378 = matrix_0_1[7] ^ matrix_0_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_380 = matrix_0_1[0] ^ _T_362; // @[AesSbox.scala 40:63]
  wire  _T_382 = matrix_0_1[1] ^ matrix_0_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_384 = _T_350 ^ _T_382; // @[AesSbox.scala 40:63]
  wire  _T_386 = _T_354 ^ _T_376; // @[AesSbox.scala 40:63]
  wire  _T_388 = _T_348 ^ _T_372; // @[AesSbox.scala 40:63]
  wire  _T_390 = matrix_0_1[7] ^ _T_354; // @[AesSbox.scala 40:63]
  wire  _T_392 = _T_388 ^ _T_356; // @[AesSbox.scala 40:63]
  wire  _T_394 = _T_388 ^ _T_360; // @[AesSbox.scala 40:63]
  wire  _T_396 = _T_360 ^ _T_384; // @[AesSbox.scala 40:63]
  wire  _T_398 = _T_378 ^ _T_374; // @[AesSbox.scala 40:63]
  wire  _T_400 = _T_390 ^ _T_380; // @[AesSbox.scala 40:63]
  wire  _T_402 = _T_384 & _T_356; // @[AesSbox.scala 41:63]
  wire  _T_404 = _T_386 & _T_368; // @[AesSbox.scala 41:63]
  wire  _T_406 = _T_370 ^ _T_402; // @[AesSbox.scala 40:63]
  wire  _T_408 = _T_366 & matrix_0_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_410 = _T_408 ^ _T_402; // @[AesSbox.scala 40:63]
  wire  _T_412 = _T_360 & _T_388; // @[AesSbox.scala 41:63]
  wire  _T_414 = _T_364 & _T_354; // @[AesSbox.scala 41:63]
  wire  _T_416 = _T_394 ^ _T_412; // @[AesSbox.scala 40:63]
  wire  _T_418 = _T_390 & _T_380; // @[AesSbox.scala 41:63]
  wire  _T_420 = _T_418 ^ _T_412; // @[AesSbox.scala 40:63]
  wire  _T_422 = _T_350 & _T_362; // @[AesSbox.scala 41:63]
  wire  _T_424 = _T_396 & _T_392; // @[AesSbox.scala 41:63]
  wire  _T_426 = _T_424 ^ _T_422; // @[AesSbox.scala 40:63]
  wire  _T_428 = _T_378 & _T_374; // @[AesSbox.scala 41:63]
  wire  _T_430 = _T_428 ^ _T_422; // @[AesSbox.scala 40:63]
  wire  _T_432 = _T_406 ^ _T_404; // @[AesSbox.scala 40:63]
  wire  _T_434 = _T_410 ^ _T_398; // @[AesSbox.scala 40:63]
  wire  _T_436 = _T_416 ^ _T_414; // @[AesSbox.scala 40:63]
  wire  _T_438 = _T_420 ^ _T_430; // @[AesSbox.scala 40:63]
  wire  _T_440 = _T_432 ^ _T_426; // @[AesSbox.scala 40:63]
  wire  _T_442 = _T_434 ^ _T_430; // @[AesSbox.scala 40:63]
  wire  _T_444 = _T_436 ^ _T_426; // @[AesSbox.scala 40:63]
  wire  _T_446 = _T_438 ^ _T_400; // @[AesSbox.scala 40:63]
  wire  _T_448 = _T_444 ^ _T_446; // @[AesSbox.scala 40:63]
  wire  _T_450 = _T_444 & _T_440; // @[AesSbox.scala 41:63]
  wire  _T_452 = _T_442 ^ _T_450; // @[AesSbox.scala 40:63]
  wire  _T_454 = _T_440 ^ _T_442; // @[AesSbox.scala 40:63]
  wire  _T_456 = _T_446 ^ _T_450; // @[AesSbox.scala 40:63]
  wire  _T_458 = _T_456 & _T_454; // @[AesSbox.scala 41:63]
  wire  _T_460 = _T_452 & _T_448; // @[AesSbox.scala 41:63]
  wire  _T_462 = _T_440 & _T_446; // @[AesSbox.scala 41:63]
  wire  _T_464 = _T_454 & _T_462; // @[AesSbox.scala 41:63]
  wire  _T_466 = _T_454 ^ _T_450; // @[AesSbox.scala 40:63]
  wire  _T_468 = _T_442 & _T_444; // @[AesSbox.scala 41:63]
  wire  _T_470 = _T_448 & _T_468; // @[AesSbox.scala 41:63]
  wire  _T_472 = _T_448 ^ _T_450; // @[AesSbox.scala 40:63]
  wire  _T_474 = _T_442 ^ _T_458; // @[AesSbox.scala 40:63]
  wire  _T_476 = _T_464 ^ _T_466; // @[AesSbox.scala 40:63]
  wire  _T_478 = _T_446 ^ _T_460; // @[AesSbox.scala 40:63]
  wire  _T_480 = _T_470 ^ _T_472; // @[AesSbox.scala 40:63]
  wire  _T_482 = _T_476 ^ _T_480; // @[AesSbox.scala 40:63]
  wire  _T_484 = _T_474 ^ _T_478; // @[AesSbox.scala 40:63]
  wire  _T_486 = _T_474 ^ _T_476; // @[AesSbox.scala 40:63]
  wire  _T_488 = _T_478 ^ _T_480; // @[AesSbox.scala 40:63]
  wire  _T_490 = _T_484 ^ _T_482; // @[AesSbox.scala 40:63]
  wire  _T_492 = _T_488 & _T_356; // @[AesSbox.scala 41:63]
  wire  _T_494 = _T_480 & _T_368; // @[AesSbox.scala 41:63]
  wire  _T_496 = _T_478 & matrix_0_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_498 = _T_486 & _T_388; // @[AesSbox.scala 41:63]
  wire  _T_500 = _T_476 & _T_354; // @[AesSbox.scala 41:63]
  wire  _T_502 = _T_474 & _T_380; // @[AesSbox.scala 41:63]
  wire  _T_504 = _T_484 & _T_362; // @[AesSbox.scala 41:63]
  wire  _T_506 = _T_490 & _T_392; // @[AesSbox.scala 41:63]
  wire  _T_508 = _T_482 & _T_374; // @[AesSbox.scala 41:63]
  wire  _T_510 = _T_488 & _T_384; // @[AesSbox.scala 41:63]
  wire  _T_512 = _T_480 & _T_386; // @[AesSbox.scala 41:63]
  wire  _T_514 = _T_478 & _T_366; // @[AesSbox.scala 41:63]
  wire  _T_516 = _T_486 & _T_360; // @[AesSbox.scala 41:63]
  wire  _T_518 = _T_476 & _T_364; // @[AesSbox.scala 41:63]
  wire  _T_520 = _T_474 & _T_390; // @[AesSbox.scala 41:63]
  wire  _T_522 = _T_484 & _T_350; // @[AesSbox.scala 41:63]
  wire  _T_524 = _T_490 & _T_396; // @[AesSbox.scala 41:63]
  wire  _T_526 = _T_482 & _T_378; // @[AesSbox.scala 41:63]
  wire  _T_528 = _T_522 ^ _T_524; // @[AesSbox.scala 40:63]
  wire  _T_530 = _T_500 ^ _T_512; // @[AesSbox.scala 40:63]
  wire  _T_532 = _T_506 ^ _T_528; // @[AesSbox.scala 40:63]
  wire  _T_534 = _T_510 ^ _T_530; // @[AesSbox.scala 40:63]
  wire  _T_536 = _T_496 ^ _T_516; // @[AesSbox.scala 40:63]
  wire  _T_538 = _T_492 ^ _T_498; // @[AesSbox.scala 40:63]
  wire  _T_540 = _T_528 ^ _T_538; // @[AesSbox.scala 40:63]
  wire  _T_542 = _T_494 ^ _T_534; // @[AesSbox.scala 40:63]
  wire  _T_544 = _T_492 ^ _T_504; // @[AesSbox.scala 40:63]
  wire  _T_546 = _T_502 ^ _T_518; // @[AesSbox.scala 40:63]
  wire  _T_548 = _T_508 ^ _T_520; // @[AesSbox.scala 40:63]
  wire  _T_550 = _T_496 ^ _T_542; // @[AesSbox.scala 40:63]
  wire  _T_552 = _T_536 ^ _T_548; // @[AesSbox.scala 40:63]
  wire  _T_554 = _T_514 ^ _T_530; // @[AesSbox.scala 40:63]
  wire  _T_556 = _T_498 ^ _T_504; // @[AesSbox.scala 40:63]
  wire  _T_558 = _T_534 ^ _T_556; // @[AesSbox.scala 40:63]
  wire  _T_560 = _T_526 ^ _T_552; // @[AesSbox.scala 40:63]
  wire  _T_562 = _T_522 ^ _T_544; // @[AesSbox.scala 40:63]
  wire  _T_564 = _T_536 ^ _T_546; // @[AesSbox.scala 40:63]
  wire  _T_565 = _T_532 ^ _T_558; // @[AesSbox.scala 40:63]
  wire  _T_566 = _T_560 ^ _T_562; // @[AesSbox.scala 42:65]
  wire  _T_567 = ~_T_566; // @[AesSbox.scala 42:51]
  wire  _T_569 = _T_502 ^ _T_528; // @[AesSbox.scala 40:63]
  wire  _T_570 = _T_540 ^ _T_542; // @[AesSbox.scala 40:63]
  wire  _T_571 = _T_550 ^ _T_569; // @[AesSbox.scala 40:63]
  wire  _T_573 = _T_500 ^ _T_516; // @[AesSbox.scala 40:63]
  wire  _T_575 = _T_538 ^ _T_554; // @[AesSbox.scala 40:63]
  wire  _T_576 = _T_540 ^ _T_564; // @[AesSbox.scala 42:65]
  wire  _T_577 = ~_T_576; // @[AesSbox.scala 42:51]
  wire  _T_579 = _T_508 ^ _T_546; // @[AesSbox.scala 40:63]
  wire  _T_581 = _T_573 ^ _T_579; // @[AesSbox.scala 40:63]
  wire  _T_583 = _T_500 ^ _T_544; // @[AesSbox.scala 40:63]
  wire  _T_584 = _T_532 ^ _T_581; // @[AesSbox.scala 42:65]
  wire  _T_585 = ~_T_584; // @[AesSbox.scala 42:51]
  wire  _T_587 = _T_552 ^ _T_575; // @[AesSbox.scala 40:63]
  wire  _T_588 = _T_532 ^ _T_587; // @[AesSbox.scala 40:63]
  wire  _T_590 = _T_542 ^ _T_583; // @[AesSbox.scala 40:63]
  wire  _T_591 = _T_532 ^ _T_590; // @[AesSbox.scala 42:65]
  wire  _T_592 = ~_T_591; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_3_1 = {_T_565,_T_592,_T_567,_T_570,_T_571,_T_588,_T_585,_T_577}; // @[Cat.scala 29:58]
  wire  _T_617 = matrix_0_2[1] ^ matrix_0_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_619 = matrix_0_2[4] ^ matrix_0_2[7]; // @[AesSbox.scala 40:63]
  wire  _T_621 = matrix_0_2[6] ^ matrix_0_2[5]; // @[AesSbox.scala 40:63]
  wire  _T_623 = matrix_0_2[0] ^ _T_621; // @[AesSbox.scala 40:63]
  wire  _T_625 = _T_617 ^ _T_619; // @[AesSbox.scala 40:63]
  wire  _T_627 = matrix_0_2[6] ^ matrix_0_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_629 = matrix_0_2[7] ^ matrix_0_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_631 = _T_617 ^ _T_627; // @[AesSbox.scala 40:63]
  wire  _T_633 = matrix_0_2[1] ^ _T_623; // @[AesSbox.scala 40:63]
  wire  _T_635 = matrix_0_2[4] ^ _T_623; // @[AesSbox.scala 40:63]
  wire  _T_637 = matrix_0_2[0] ^ _T_625; // @[AesSbox.scala 40:63]
  wire  _T_639 = _T_625 ^ _T_627; // @[AesSbox.scala 40:63]
  wire  _T_641 = matrix_0_2[5] ^ matrix_0_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_643 = _T_621 ^ _T_625; // @[AesSbox.scala 40:63]
  wire  _T_645 = matrix_0_2[2] ^ _T_629; // @[AesSbox.scala 40:63]
  wire  _T_647 = matrix_0_2[7] ^ matrix_0_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_649 = matrix_0_2[0] ^ _T_631; // @[AesSbox.scala 40:63]
  wire  _T_651 = matrix_0_2[1] ^ matrix_0_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_653 = _T_619 ^ _T_651; // @[AesSbox.scala 40:63]
  wire  _T_655 = _T_623 ^ _T_645; // @[AesSbox.scala 40:63]
  wire  _T_657 = _T_617 ^ _T_641; // @[AesSbox.scala 40:63]
  wire  _T_659 = matrix_0_2[7] ^ _T_623; // @[AesSbox.scala 40:63]
  wire  _T_661 = _T_657 ^ _T_625; // @[AesSbox.scala 40:63]
  wire  _T_663 = _T_657 ^ _T_629; // @[AesSbox.scala 40:63]
  wire  _T_665 = _T_629 ^ _T_653; // @[AesSbox.scala 40:63]
  wire  _T_667 = _T_647 ^ _T_643; // @[AesSbox.scala 40:63]
  wire  _T_669 = _T_659 ^ _T_649; // @[AesSbox.scala 40:63]
  wire  _T_671 = _T_653 & _T_625; // @[AesSbox.scala 41:63]
  wire  _T_673 = _T_655 & _T_637; // @[AesSbox.scala 41:63]
  wire  _T_675 = _T_639 ^ _T_671; // @[AesSbox.scala 40:63]
  wire  _T_677 = _T_635 & matrix_0_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_679 = _T_677 ^ _T_671; // @[AesSbox.scala 40:63]
  wire  _T_681 = _T_629 & _T_657; // @[AesSbox.scala 41:63]
  wire  _T_683 = _T_633 & _T_623; // @[AesSbox.scala 41:63]
  wire  _T_685 = _T_663 ^ _T_681; // @[AesSbox.scala 40:63]
  wire  _T_687 = _T_659 & _T_649; // @[AesSbox.scala 41:63]
  wire  _T_689 = _T_687 ^ _T_681; // @[AesSbox.scala 40:63]
  wire  _T_691 = _T_619 & _T_631; // @[AesSbox.scala 41:63]
  wire  _T_693 = _T_665 & _T_661; // @[AesSbox.scala 41:63]
  wire  _T_695 = _T_693 ^ _T_691; // @[AesSbox.scala 40:63]
  wire  _T_697 = _T_647 & _T_643; // @[AesSbox.scala 41:63]
  wire  _T_699 = _T_697 ^ _T_691; // @[AesSbox.scala 40:63]
  wire  _T_701 = _T_675 ^ _T_673; // @[AesSbox.scala 40:63]
  wire  _T_703 = _T_679 ^ _T_667; // @[AesSbox.scala 40:63]
  wire  _T_705 = _T_685 ^ _T_683; // @[AesSbox.scala 40:63]
  wire  _T_707 = _T_689 ^ _T_699; // @[AesSbox.scala 40:63]
  wire  _T_709 = _T_701 ^ _T_695; // @[AesSbox.scala 40:63]
  wire  _T_711 = _T_703 ^ _T_699; // @[AesSbox.scala 40:63]
  wire  _T_713 = _T_705 ^ _T_695; // @[AesSbox.scala 40:63]
  wire  _T_715 = _T_707 ^ _T_669; // @[AesSbox.scala 40:63]
  wire  _T_717 = _T_713 ^ _T_715; // @[AesSbox.scala 40:63]
  wire  _T_719 = _T_713 & _T_709; // @[AesSbox.scala 41:63]
  wire  _T_721 = _T_711 ^ _T_719; // @[AesSbox.scala 40:63]
  wire  _T_723 = _T_709 ^ _T_711; // @[AesSbox.scala 40:63]
  wire  _T_725 = _T_715 ^ _T_719; // @[AesSbox.scala 40:63]
  wire  _T_727 = _T_725 & _T_723; // @[AesSbox.scala 41:63]
  wire  _T_729 = _T_721 & _T_717; // @[AesSbox.scala 41:63]
  wire  _T_731 = _T_709 & _T_715; // @[AesSbox.scala 41:63]
  wire  _T_733 = _T_723 & _T_731; // @[AesSbox.scala 41:63]
  wire  _T_735 = _T_723 ^ _T_719; // @[AesSbox.scala 40:63]
  wire  _T_737 = _T_711 & _T_713; // @[AesSbox.scala 41:63]
  wire  _T_739 = _T_717 & _T_737; // @[AesSbox.scala 41:63]
  wire  _T_741 = _T_717 ^ _T_719; // @[AesSbox.scala 40:63]
  wire  _T_743 = _T_711 ^ _T_727; // @[AesSbox.scala 40:63]
  wire  _T_745 = _T_733 ^ _T_735; // @[AesSbox.scala 40:63]
  wire  _T_747 = _T_715 ^ _T_729; // @[AesSbox.scala 40:63]
  wire  _T_749 = _T_739 ^ _T_741; // @[AesSbox.scala 40:63]
  wire  _T_751 = _T_745 ^ _T_749; // @[AesSbox.scala 40:63]
  wire  _T_753 = _T_743 ^ _T_747; // @[AesSbox.scala 40:63]
  wire  _T_755 = _T_743 ^ _T_745; // @[AesSbox.scala 40:63]
  wire  _T_757 = _T_747 ^ _T_749; // @[AesSbox.scala 40:63]
  wire  _T_759 = _T_753 ^ _T_751; // @[AesSbox.scala 40:63]
  wire  _T_761 = _T_757 & _T_625; // @[AesSbox.scala 41:63]
  wire  _T_763 = _T_749 & _T_637; // @[AesSbox.scala 41:63]
  wire  _T_765 = _T_747 & matrix_0_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_767 = _T_755 & _T_657; // @[AesSbox.scala 41:63]
  wire  _T_769 = _T_745 & _T_623; // @[AesSbox.scala 41:63]
  wire  _T_771 = _T_743 & _T_649; // @[AesSbox.scala 41:63]
  wire  _T_773 = _T_753 & _T_631; // @[AesSbox.scala 41:63]
  wire  _T_775 = _T_759 & _T_661; // @[AesSbox.scala 41:63]
  wire  _T_777 = _T_751 & _T_643; // @[AesSbox.scala 41:63]
  wire  _T_779 = _T_757 & _T_653; // @[AesSbox.scala 41:63]
  wire  _T_781 = _T_749 & _T_655; // @[AesSbox.scala 41:63]
  wire  _T_783 = _T_747 & _T_635; // @[AesSbox.scala 41:63]
  wire  _T_785 = _T_755 & _T_629; // @[AesSbox.scala 41:63]
  wire  _T_787 = _T_745 & _T_633; // @[AesSbox.scala 41:63]
  wire  _T_789 = _T_743 & _T_659; // @[AesSbox.scala 41:63]
  wire  _T_791 = _T_753 & _T_619; // @[AesSbox.scala 41:63]
  wire  _T_793 = _T_759 & _T_665; // @[AesSbox.scala 41:63]
  wire  _T_795 = _T_751 & _T_647; // @[AesSbox.scala 41:63]
  wire  _T_797 = _T_791 ^ _T_793; // @[AesSbox.scala 40:63]
  wire  _T_799 = _T_769 ^ _T_781; // @[AesSbox.scala 40:63]
  wire  _T_801 = _T_775 ^ _T_797; // @[AesSbox.scala 40:63]
  wire  _T_803 = _T_779 ^ _T_799; // @[AesSbox.scala 40:63]
  wire  _T_805 = _T_765 ^ _T_785; // @[AesSbox.scala 40:63]
  wire  _T_807 = _T_761 ^ _T_767; // @[AesSbox.scala 40:63]
  wire  _T_809 = _T_797 ^ _T_807; // @[AesSbox.scala 40:63]
  wire  _T_811 = _T_763 ^ _T_803; // @[AesSbox.scala 40:63]
  wire  _T_813 = _T_761 ^ _T_773; // @[AesSbox.scala 40:63]
  wire  _T_815 = _T_771 ^ _T_787; // @[AesSbox.scala 40:63]
  wire  _T_817 = _T_777 ^ _T_789; // @[AesSbox.scala 40:63]
  wire  _T_819 = _T_765 ^ _T_811; // @[AesSbox.scala 40:63]
  wire  _T_821 = _T_805 ^ _T_817; // @[AesSbox.scala 40:63]
  wire  _T_823 = _T_783 ^ _T_799; // @[AesSbox.scala 40:63]
  wire  _T_825 = _T_767 ^ _T_773; // @[AesSbox.scala 40:63]
  wire  _T_827 = _T_803 ^ _T_825; // @[AesSbox.scala 40:63]
  wire  _T_829 = _T_795 ^ _T_821; // @[AesSbox.scala 40:63]
  wire  _T_831 = _T_791 ^ _T_813; // @[AesSbox.scala 40:63]
  wire  _T_833 = _T_805 ^ _T_815; // @[AesSbox.scala 40:63]
  wire  _T_834 = _T_801 ^ _T_827; // @[AesSbox.scala 40:63]
  wire  _T_835 = _T_829 ^ _T_831; // @[AesSbox.scala 42:65]
  wire  _T_836 = ~_T_835; // @[AesSbox.scala 42:51]
  wire  _T_838 = _T_771 ^ _T_797; // @[AesSbox.scala 40:63]
  wire  _T_839 = _T_809 ^ _T_811; // @[AesSbox.scala 40:63]
  wire  _T_840 = _T_819 ^ _T_838; // @[AesSbox.scala 40:63]
  wire  _T_842 = _T_769 ^ _T_785; // @[AesSbox.scala 40:63]
  wire  _T_844 = _T_807 ^ _T_823; // @[AesSbox.scala 40:63]
  wire  _T_845 = _T_809 ^ _T_833; // @[AesSbox.scala 42:65]
  wire  _T_846 = ~_T_845; // @[AesSbox.scala 42:51]
  wire  _T_848 = _T_777 ^ _T_815; // @[AesSbox.scala 40:63]
  wire  _T_850 = _T_842 ^ _T_848; // @[AesSbox.scala 40:63]
  wire  _T_852 = _T_769 ^ _T_813; // @[AesSbox.scala 40:63]
  wire  _T_853 = _T_801 ^ _T_850; // @[AesSbox.scala 42:65]
  wire  _T_854 = ~_T_853; // @[AesSbox.scala 42:51]
  wire  _T_856 = _T_821 ^ _T_844; // @[AesSbox.scala 40:63]
  wire  _T_857 = _T_801 ^ _T_856; // @[AesSbox.scala 40:63]
  wire  _T_859 = _T_811 ^ _T_852; // @[AesSbox.scala 40:63]
  wire  _T_860 = _T_801 ^ _T_859; // @[AesSbox.scala 42:65]
  wire  _T_861 = ~_T_860; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_2_2 = {_T_834,_T_861,_T_836,_T_839,_T_840,_T_857,_T_854,_T_846}; // @[Cat.scala 29:58]
  wire  _T_886 = matrix_0_3[1] ^ matrix_0_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_888 = matrix_0_3[4] ^ matrix_0_3[7]; // @[AesSbox.scala 40:63]
  wire  _T_890 = matrix_0_3[6] ^ matrix_0_3[5]; // @[AesSbox.scala 40:63]
  wire  _T_892 = matrix_0_3[0] ^ _T_890; // @[AesSbox.scala 40:63]
  wire  _T_894 = _T_886 ^ _T_888; // @[AesSbox.scala 40:63]
  wire  _T_896 = matrix_0_3[6] ^ matrix_0_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_898 = matrix_0_3[7] ^ matrix_0_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_900 = _T_886 ^ _T_896; // @[AesSbox.scala 40:63]
  wire  _T_902 = matrix_0_3[1] ^ _T_892; // @[AesSbox.scala 40:63]
  wire  _T_904 = matrix_0_3[4] ^ _T_892; // @[AesSbox.scala 40:63]
  wire  _T_906 = matrix_0_3[0] ^ _T_894; // @[AesSbox.scala 40:63]
  wire  _T_908 = _T_894 ^ _T_896; // @[AesSbox.scala 40:63]
  wire  _T_910 = matrix_0_3[5] ^ matrix_0_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_912 = _T_890 ^ _T_894; // @[AesSbox.scala 40:63]
  wire  _T_914 = matrix_0_3[2] ^ _T_898; // @[AesSbox.scala 40:63]
  wire  _T_916 = matrix_0_3[7] ^ matrix_0_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_918 = matrix_0_3[0] ^ _T_900; // @[AesSbox.scala 40:63]
  wire  _T_920 = matrix_0_3[1] ^ matrix_0_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_922 = _T_888 ^ _T_920; // @[AesSbox.scala 40:63]
  wire  _T_924 = _T_892 ^ _T_914; // @[AesSbox.scala 40:63]
  wire  _T_926 = _T_886 ^ _T_910; // @[AesSbox.scala 40:63]
  wire  _T_928 = matrix_0_3[7] ^ _T_892; // @[AesSbox.scala 40:63]
  wire  _T_930 = _T_926 ^ _T_894; // @[AesSbox.scala 40:63]
  wire  _T_932 = _T_926 ^ _T_898; // @[AesSbox.scala 40:63]
  wire  _T_934 = _T_898 ^ _T_922; // @[AesSbox.scala 40:63]
  wire  _T_936 = _T_916 ^ _T_912; // @[AesSbox.scala 40:63]
  wire  _T_938 = _T_928 ^ _T_918; // @[AesSbox.scala 40:63]
  wire  _T_940 = _T_922 & _T_894; // @[AesSbox.scala 41:63]
  wire  _T_942 = _T_924 & _T_906; // @[AesSbox.scala 41:63]
  wire  _T_944 = _T_908 ^ _T_940; // @[AesSbox.scala 40:63]
  wire  _T_946 = _T_904 & matrix_0_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_948 = _T_946 ^ _T_940; // @[AesSbox.scala 40:63]
  wire  _T_950 = _T_898 & _T_926; // @[AesSbox.scala 41:63]
  wire  _T_952 = _T_902 & _T_892; // @[AesSbox.scala 41:63]
  wire  _T_954 = _T_932 ^ _T_950; // @[AesSbox.scala 40:63]
  wire  _T_956 = _T_928 & _T_918; // @[AesSbox.scala 41:63]
  wire  _T_958 = _T_956 ^ _T_950; // @[AesSbox.scala 40:63]
  wire  _T_960 = _T_888 & _T_900; // @[AesSbox.scala 41:63]
  wire  _T_962 = _T_934 & _T_930; // @[AesSbox.scala 41:63]
  wire  _T_964 = _T_962 ^ _T_960; // @[AesSbox.scala 40:63]
  wire  _T_966 = _T_916 & _T_912; // @[AesSbox.scala 41:63]
  wire  _T_968 = _T_966 ^ _T_960; // @[AesSbox.scala 40:63]
  wire  _T_970 = _T_944 ^ _T_942; // @[AesSbox.scala 40:63]
  wire  _T_972 = _T_948 ^ _T_936; // @[AesSbox.scala 40:63]
  wire  _T_974 = _T_954 ^ _T_952; // @[AesSbox.scala 40:63]
  wire  _T_976 = _T_958 ^ _T_968; // @[AesSbox.scala 40:63]
  wire  _T_978 = _T_970 ^ _T_964; // @[AesSbox.scala 40:63]
  wire  _T_980 = _T_972 ^ _T_968; // @[AesSbox.scala 40:63]
  wire  _T_982 = _T_974 ^ _T_964; // @[AesSbox.scala 40:63]
  wire  _T_984 = _T_976 ^ _T_938; // @[AesSbox.scala 40:63]
  wire  _T_986 = _T_982 ^ _T_984; // @[AesSbox.scala 40:63]
  wire  _T_988 = _T_982 & _T_978; // @[AesSbox.scala 41:63]
  wire  _T_990 = _T_980 ^ _T_988; // @[AesSbox.scala 40:63]
  wire  _T_992 = _T_978 ^ _T_980; // @[AesSbox.scala 40:63]
  wire  _T_994 = _T_984 ^ _T_988; // @[AesSbox.scala 40:63]
  wire  _T_996 = _T_994 & _T_992; // @[AesSbox.scala 41:63]
  wire  _T_998 = _T_990 & _T_986; // @[AesSbox.scala 41:63]
  wire  _T_1000 = _T_978 & _T_984; // @[AesSbox.scala 41:63]
  wire  _T_1002 = _T_992 & _T_1000; // @[AesSbox.scala 41:63]
  wire  _T_1004 = _T_992 ^ _T_988; // @[AesSbox.scala 40:63]
  wire  _T_1006 = _T_980 & _T_982; // @[AesSbox.scala 41:63]
  wire  _T_1008 = _T_986 & _T_1006; // @[AesSbox.scala 41:63]
  wire  _T_1010 = _T_986 ^ _T_988; // @[AesSbox.scala 40:63]
  wire  _T_1012 = _T_980 ^ _T_996; // @[AesSbox.scala 40:63]
  wire  _T_1014 = _T_1002 ^ _T_1004; // @[AesSbox.scala 40:63]
  wire  _T_1016 = _T_984 ^ _T_998; // @[AesSbox.scala 40:63]
  wire  _T_1018 = _T_1008 ^ _T_1010; // @[AesSbox.scala 40:63]
  wire  _T_1020 = _T_1014 ^ _T_1018; // @[AesSbox.scala 40:63]
  wire  _T_1022 = _T_1012 ^ _T_1016; // @[AesSbox.scala 40:63]
  wire  _T_1024 = _T_1012 ^ _T_1014; // @[AesSbox.scala 40:63]
  wire  _T_1026 = _T_1016 ^ _T_1018; // @[AesSbox.scala 40:63]
  wire  _T_1028 = _T_1022 ^ _T_1020; // @[AesSbox.scala 40:63]
  wire  _T_1030 = _T_1026 & _T_894; // @[AesSbox.scala 41:63]
  wire  _T_1032 = _T_1018 & _T_906; // @[AesSbox.scala 41:63]
  wire  _T_1034 = _T_1016 & matrix_0_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_1036 = _T_1024 & _T_926; // @[AesSbox.scala 41:63]
  wire  _T_1038 = _T_1014 & _T_892; // @[AesSbox.scala 41:63]
  wire  _T_1040 = _T_1012 & _T_918; // @[AesSbox.scala 41:63]
  wire  _T_1042 = _T_1022 & _T_900; // @[AesSbox.scala 41:63]
  wire  _T_1044 = _T_1028 & _T_930; // @[AesSbox.scala 41:63]
  wire  _T_1046 = _T_1020 & _T_912; // @[AesSbox.scala 41:63]
  wire  _T_1048 = _T_1026 & _T_922; // @[AesSbox.scala 41:63]
  wire  _T_1050 = _T_1018 & _T_924; // @[AesSbox.scala 41:63]
  wire  _T_1052 = _T_1016 & _T_904; // @[AesSbox.scala 41:63]
  wire  _T_1054 = _T_1024 & _T_898; // @[AesSbox.scala 41:63]
  wire  _T_1056 = _T_1014 & _T_902; // @[AesSbox.scala 41:63]
  wire  _T_1058 = _T_1012 & _T_928; // @[AesSbox.scala 41:63]
  wire  _T_1060 = _T_1022 & _T_888; // @[AesSbox.scala 41:63]
  wire  _T_1062 = _T_1028 & _T_934; // @[AesSbox.scala 41:63]
  wire  _T_1064 = _T_1020 & _T_916; // @[AesSbox.scala 41:63]
  wire  _T_1066 = _T_1060 ^ _T_1062; // @[AesSbox.scala 40:63]
  wire  _T_1068 = _T_1038 ^ _T_1050; // @[AesSbox.scala 40:63]
  wire  _T_1070 = _T_1044 ^ _T_1066; // @[AesSbox.scala 40:63]
  wire  _T_1072 = _T_1048 ^ _T_1068; // @[AesSbox.scala 40:63]
  wire  _T_1074 = _T_1034 ^ _T_1054; // @[AesSbox.scala 40:63]
  wire  _T_1076 = _T_1030 ^ _T_1036; // @[AesSbox.scala 40:63]
  wire  _T_1078 = _T_1066 ^ _T_1076; // @[AesSbox.scala 40:63]
  wire  _T_1080 = _T_1032 ^ _T_1072; // @[AesSbox.scala 40:63]
  wire  _T_1082 = _T_1030 ^ _T_1042; // @[AesSbox.scala 40:63]
  wire  _T_1084 = _T_1040 ^ _T_1056; // @[AesSbox.scala 40:63]
  wire  _T_1086 = _T_1046 ^ _T_1058; // @[AesSbox.scala 40:63]
  wire  _T_1088 = _T_1034 ^ _T_1080; // @[AesSbox.scala 40:63]
  wire  _T_1090 = _T_1074 ^ _T_1086; // @[AesSbox.scala 40:63]
  wire  _T_1092 = _T_1052 ^ _T_1068; // @[AesSbox.scala 40:63]
  wire  _T_1094 = _T_1036 ^ _T_1042; // @[AesSbox.scala 40:63]
  wire  _T_1096 = _T_1072 ^ _T_1094; // @[AesSbox.scala 40:63]
  wire  _T_1098 = _T_1064 ^ _T_1090; // @[AesSbox.scala 40:63]
  wire  _T_1100 = _T_1060 ^ _T_1082; // @[AesSbox.scala 40:63]
  wire  _T_1102 = _T_1074 ^ _T_1084; // @[AesSbox.scala 40:63]
  wire  _T_1103 = _T_1070 ^ _T_1096; // @[AesSbox.scala 40:63]
  wire  _T_1104 = _T_1098 ^ _T_1100; // @[AesSbox.scala 42:65]
  wire  _T_1105 = ~_T_1104; // @[AesSbox.scala 42:51]
  wire  _T_1107 = _T_1040 ^ _T_1066; // @[AesSbox.scala 40:63]
  wire  _T_1108 = _T_1078 ^ _T_1080; // @[AesSbox.scala 40:63]
  wire  _T_1109 = _T_1088 ^ _T_1107; // @[AesSbox.scala 40:63]
  wire  _T_1111 = _T_1038 ^ _T_1054; // @[AesSbox.scala 40:63]
  wire  _T_1113 = _T_1076 ^ _T_1092; // @[AesSbox.scala 40:63]
  wire  _T_1114 = _T_1078 ^ _T_1102; // @[AesSbox.scala 42:65]
  wire  _T_1115 = ~_T_1114; // @[AesSbox.scala 42:51]
  wire  _T_1117 = _T_1046 ^ _T_1084; // @[AesSbox.scala 40:63]
  wire  _T_1119 = _T_1111 ^ _T_1117; // @[AesSbox.scala 40:63]
  wire  _T_1121 = _T_1038 ^ _T_1082; // @[AesSbox.scala 40:63]
  wire  _T_1122 = _T_1070 ^ _T_1119; // @[AesSbox.scala 42:65]
  wire  _T_1123 = ~_T_1122; // @[AesSbox.scala 42:51]
  wire  _T_1125 = _T_1090 ^ _T_1113; // @[AesSbox.scala 40:63]
  wire  _T_1126 = _T_1070 ^ _T_1125; // @[AesSbox.scala 40:63]
  wire  _T_1128 = _T_1080 ^ _T_1121; // @[AesSbox.scala 40:63]
  wire  _T_1129 = _T_1070 ^ _T_1128; // @[AesSbox.scala 42:65]
  wire  _T_1130 = ~_T_1129; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_1_3 = {_T_1103,_T_1130,_T_1105,_T_1108,_T_1109,_T_1126,_T_1123,_T_1115}; // @[Cat.scala 29:58]
  wire  _T_1156 = matrix_1_0[1] ^ matrix_1_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_1158 = matrix_1_0[4] ^ matrix_1_0[7]; // @[AesSbox.scala 40:63]
  wire  _T_1160 = matrix_1_0[6] ^ matrix_1_0[5]; // @[AesSbox.scala 40:63]
  wire  _T_1162 = matrix_1_0[0] ^ _T_1160; // @[AesSbox.scala 40:63]
  wire  _T_1164 = _T_1156 ^ _T_1158; // @[AesSbox.scala 40:63]
  wire  _T_1166 = matrix_1_0[6] ^ matrix_1_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_1168 = matrix_1_0[7] ^ matrix_1_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_1170 = _T_1156 ^ _T_1166; // @[AesSbox.scala 40:63]
  wire  _T_1172 = matrix_1_0[1] ^ _T_1162; // @[AesSbox.scala 40:63]
  wire  _T_1174 = matrix_1_0[4] ^ _T_1162; // @[AesSbox.scala 40:63]
  wire  _T_1176 = matrix_1_0[0] ^ _T_1164; // @[AesSbox.scala 40:63]
  wire  _T_1178 = _T_1164 ^ _T_1166; // @[AesSbox.scala 40:63]
  wire  _T_1180 = matrix_1_0[5] ^ matrix_1_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_1182 = _T_1160 ^ _T_1164; // @[AesSbox.scala 40:63]
  wire  _T_1184 = matrix_1_0[2] ^ _T_1168; // @[AesSbox.scala 40:63]
  wire  _T_1186 = matrix_1_0[7] ^ matrix_1_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_1188 = matrix_1_0[0] ^ _T_1170; // @[AesSbox.scala 40:63]
  wire  _T_1190 = matrix_1_0[1] ^ matrix_1_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_1192 = _T_1158 ^ _T_1190; // @[AesSbox.scala 40:63]
  wire  _T_1194 = _T_1162 ^ _T_1184; // @[AesSbox.scala 40:63]
  wire  _T_1196 = _T_1156 ^ _T_1180; // @[AesSbox.scala 40:63]
  wire  _T_1198 = matrix_1_0[7] ^ _T_1162; // @[AesSbox.scala 40:63]
  wire  _T_1200 = _T_1196 ^ _T_1164; // @[AesSbox.scala 40:63]
  wire  _T_1202 = _T_1196 ^ _T_1168; // @[AesSbox.scala 40:63]
  wire  _T_1204 = _T_1168 ^ _T_1192; // @[AesSbox.scala 40:63]
  wire  _T_1206 = _T_1186 ^ _T_1182; // @[AesSbox.scala 40:63]
  wire  _T_1208 = _T_1198 ^ _T_1188; // @[AesSbox.scala 40:63]
  wire  _T_1210 = _T_1192 & _T_1164; // @[AesSbox.scala 41:63]
  wire  _T_1212 = _T_1194 & _T_1176; // @[AesSbox.scala 41:63]
  wire  _T_1214 = _T_1178 ^ _T_1210; // @[AesSbox.scala 40:63]
  wire  _T_1216 = _T_1174 & matrix_1_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_1218 = _T_1216 ^ _T_1210; // @[AesSbox.scala 40:63]
  wire  _T_1220 = _T_1168 & _T_1196; // @[AesSbox.scala 41:63]
  wire  _T_1222 = _T_1172 & _T_1162; // @[AesSbox.scala 41:63]
  wire  _T_1224 = _T_1202 ^ _T_1220; // @[AesSbox.scala 40:63]
  wire  _T_1226 = _T_1198 & _T_1188; // @[AesSbox.scala 41:63]
  wire  _T_1228 = _T_1226 ^ _T_1220; // @[AesSbox.scala 40:63]
  wire  _T_1230 = _T_1158 & _T_1170; // @[AesSbox.scala 41:63]
  wire  _T_1232 = _T_1204 & _T_1200; // @[AesSbox.scala 41:63]
  wire  _T_1234 = _T_1232 ^ _T_1230; // @[AesSbox.scala 40:63]
  wire  _T_1236 = _T_1186 & _T_1182; // @[AesSbox.scala 41:63]
  wire  _T_1238 = _T_1236 ^ _T_1230; // @[AesSbox.scala 40:63]
  wire  _T_1240 = _T_1214 ^ _T_1212; // @[AesSbox.scala 40:63]
  wire  _T_1242 = _T_1218 ^ _T_1206; // @[AesSbox.scala 40:63]
  wire  _T_1244 = _T_1224 ^ _T_1222; // @[AesSbox.scala 40:63]
  wire  _T_1246 = _T_1228 ^ _T_1238; // @[AesSbox.scala 40:63]
  wire  _T_1248 = _T_1240 ^ _T_1234; // @[AesSbox.scala 40:63]
  wire  _T_1250 = _T_1242 ^ _T_1238; // @[AesSbox.scala 40:63]
  wire  _T_1252 = _T_1244 ^ _T_1234; // @[AesSbox.scala 40:63]
  wire  _T_1254 = _T_1246 ^ _T_1208; // @[AesSbox.scala 40:63]
  wire  _T_1256 = _T_1252 ^ _T_1254; // @[AesSbox.scala 40:63]
  wire  _T_1258 = _T_1252 & _T_1248; // @[AesSbox.scala 41:63]
  wire  _T_1260 = _T_1250 ^ _T_1258; // @[AesSbox.scala 40:63]
  wire  _T_1262 = _T_1248 ^ _T_1250; // @[AesSbox.scala 40:63]
  wire  _T_1264 = _T_1254 ^ _T_1258; // @[AesSbox.scala 40:63]
  wire  _T_1266 = _T_1264 & _T_1262; // @[AesSbox.scala 41:63]
  wire  _T_1268 = _T_1260 & _T_1256; // @[AesSbox.scala 41:63]
  wire  _T_1270 = _T_1248 & _T_1254; // @[AesSbox.scala 41:63]
  wire  _T_1272 = _T_1262 & _T_1270; // @[AesSbox.scala 41:63]
  wire  _T_1274 = _T_1262 ^ _T_1258; // @[AesSbox.scala 40:63]
  wire  _T_1276 = _T_1250 & _T_1252; // @[AesSbox.scala 41:63]
  wire  _T_1278 = _T_1256 & _T_1276; // @[AesSbox.scala 41:63]
  wire  _T_1280 = _T_1256 ^ _T_1258; // @[AesSbox.scala 40:63]
  wire  _T_1282 = _T_1250 ^ _T_1266; // @[AesSbox.scala 40:63]
  wire  _T_1284 = _T_1272 ^ _T_1274; // @[AesSbox.scala 40:63]
  wire  _T_1286 = _T_1254 ^ _T_1268; // @[AesSbox.scala 40:63]
  wire  _T_1288 = _T_1278 ^ _T_1280; // @[AesSbox.scala 40:63]
  wire  _T_1290 = _T_1284 ^ _T_1288; // @[AesSbox.scala 40:63]
  wire  _T_1292 = _T_1282 ^ _T_1286; // @[AesSbox.scala 40:63]
  wire  _T_1294 = _T_1282 ^ _T_1284; // @[AesSbox.scala 40:63]
  wire  _T_1296 = _T_1286 ^ _T_1288; // @[AesSbox.scala 40:63]
  wire  _T_1298 = _T_1292 ^ _T_1290; // @[AesSbox.scala 40:63]
  wire  _T_1300 = _T_1296 & _T_1164; // @[AesSbox.scala 41:63]
  wire  _T_1302 = _T_1288 & _T_1176; // @[AesSbox.scala 41:63]
  wire  _T_1304 = _T_1286 & matrix_1_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_1306 = _T_1294 & _T_1196; // @[AesSbox.scala 41:63]
  wire  _T_1308 = _T_1284 & _T_1162; // @[AesSbox.scala 41:63]
  wire  _T_1310 = _T_1282 & _T_1188; // @[AesSbox.scala 41:63]
  wire  _T_1312 = _T_1292 & _T_1170; // @[AesSbox.scala 41:63]
  wire  _T_1314 = _T_1298 & _T_1200; // @[AesSbox.scala 41:63]
  wire  _T_1316 = _T_1290 & _T_1182; // @[AesSbox.scala 41:63]
  wire  _T_1318 = _T_1296 & _T_1192; // @[AesSbox.scala 41:63]
  wire  _T_1320 = _T_1288 & _T_1194; // @[AesSbox.scala 41:63]
  wire  _T_1322 = _T_1286 & _T_1174; // @[AesSbox.scala 41:63]
  wire  _T_1324 = _T_1294 & _T_1168; // @[AesSbox.scala 41:63]
  wire  _T_1326 = _T_1284 & _T_1172; // @[AesSbox.scala 41:63]
  wire  _T_1328 = _T_1282 & _T_1198; // @[AesSbox.scala 41:63]
  wire  _T_1330 = _T_1292 & _T_1158; // @[AesSbox.scala 41:63]
  wire  _T_1332 = _T_1298 & _T_1204; // @[AesSbox.scala 41:63]
  wire  _T_1334 = _T_1290 & _T_1186; // @[AesSbox.scala 41:63]
  wire  _T_1336 = _T_1330 ^ _T_1332; // @[AesSbox.scala 40:63]
  wire  _T_1338 = _T_1308 ^ _T_1320; // @[AesSbox.scala 40:63]
  wire  _T_1340 = _T_1314 ^ _T_1336; // @[AesSbox.scala 40:63]
  wire  _T_1342 = _T_1318 ^ _T_1338; // @[AesSbox.scala 40:63]
  wire  _T_1344 = _T_1304 ^ _T_1324; // @[AesSbox.scala 40:63]
  wire  _T_1346 = _T_1300 ^ _T_1306; // @[AesSbox.scala 40:63]
  wire  _T_1348 = _T_1336 ^ _T_1346; // @[AesSbox.scala 40:63]
  wire  _T_1350 = _T_1302 ^ _T_1342; // @[AesSbox.scala 40:63]
  wire  _T_1352 = _T_1300 ^ _T_1312; // @[AesSbox.scala 40:63]
  wire  _T_1354 = _T_1310 ^ _T_1326; // @[AesSbox.scala 40:63]
  wire  _T_1356 = _T_1316 ^ _T_1328; // @[AesSbox.scala 40:63]
  wire  _T_1358 = _T_1304 ^ _T_1350; // @[AesSbox.scala 40:63]
  wire  _T_1360 = _T_1344 ^ _T_1356; // @[AesSbox.scala 40:63]
  wire  _T_1362 = _T_1322 ^ _T_1338; // @[AesSbox.scala 40:63]
  wire  _T_1364 = _T_1306 ^ _T_1312; // @[AesSbox.scala 40:63]
  wire  _T_1366 = _T_1342 ^ _T_1364; // @[AesSbox.scala 40:63]
  wire  _T_1368 = _T_1334 ^ _T_1360; // @[AesSbox.scala 40:63]
  wire  _T_1370 = _T_1330 ^ _T_1352; // @[AesSbox.scala 40:63]
  wire  _T_1372 = _T_1344 ^ _T_1354; // @[AesSbox.scala 40:63]
  wire  _T_1373 = _T_1340 ^ _T_1366; // @[AesSbox.scala 40:63]
  wire  _T_1374 = _T_1368 ^ _T_1370; // @[AesSbox.scala 42:65]
  wire  _T_1375 = ~_T_1374; // @[AesSbox.scala 42:51]
  wire  _T_1377 = _T_1310 ^ _T_1336; // @[AesSbox.scala 40:63]
  wire  _T_1378 = _T_1348 ^ _T_1350; // @[AesSbox.scala 40:63]
  wire  _T_1379 = _T_1358 ^ _T_1377; // @[AesSbox.scala 40:63]
  wire  _T_1381 = _T_1308 ^ _T_1324; // @[AesSbox.scala 40:63]
  wire  _T_1383 = _T_1346 ^ _T_1362; // @[AesSbox.scala 40:63]
  wire  _T_1384 = _T_1348 ^ _T_1372; // @[AesSbox.scala 42:65]
  wire  _T_1385 = ~_T_1384; // @[AesSbox.scala 42:51]
  wire  _T_1387 = _T_1316 ^ _T_1354; // @[AesSbox.scala 40:63]
  wire  _T_1389 = _T_1381 ^ _T_1387; // @[AesSbox.scala 40:63]
  wire  _T_1391 = _T_1308 ^ _T_1352; // @[AesSbox.scala 40:63]
  wire  _T_1392 = _T_1340 ^ _T_1389; // @[AesSbox.scala 42:65]
  wire  _T_1393 = ~_T_1392; // @[AesSbox.scala 42:51]
  wire  _T_1395 = _T_1360 ^ _T_1383; // @[AesSbox.scala 40:63]
  wire  _T_1396 = _T_1340 ^ _T_1395; // @[AesSbox.scala 40:63]
  wire  _T_1398 = _T_1350 ^ _T_1391; // @[AesSbox.scala 40:63]
  wire  _T_1399 = _T_1340 ^ _T_1398; // @[AesSbox.scala 42:65]
  wire  _T_1400 = ~_T_1399; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_1_0 = {_T_1373,_T_1400,_T_1375,_T_1378,_T_1379,_T_1396,_T_1393,_T_1385}; // @[Cat.scala 29:58]
  wire  _T_1425 = matrix_1_1[1] ^ matrix_1_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_1427 = matrix_1_1[4] ^ matrix_1_1[7]; // @[AesSbox.scala 40:63]
  wire  _T_1429 = matrix_1_1[6] ^ matrix_1_1[5]; // @[AesSbox.scala 40:63]
  wire  _T_1431 = matrix_1_1[0] ^ _T_1429; // @[AesSbox.scala 40:63]
  wire  _T_1433 = _T_1425 ^ _T_1427; // @[AesSbox.scala 40:63]
  wire  _T_1435 = matrix_1_1[6] ^ matrix_1_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_1437 = matrix_1_1[7] ^ matrix_1_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_1439 = _T_1425 ^ _T_1435; // @[AesSbox.scala 40:63]
  wire  _T_1441 = matrix_1_1[1] ^ _T_1431; // @[AesSbox.scala 40:63]
  wire  _T_1443 = matrix_1_1[4] ^ _T_1431; // @[AesSbox.scala 40:63]
  wire  _T_1445 = matrix_1_1[0] ^ _T_1433; // @[AesSbox.scala 40:63]
  wire  _T_1447 = _T_1433 ^ _T_1435; // @[AesSbox.scala 40:63]
  wire  _T_1449 = matrix_1_1[5] ^ matrix_1_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_1451 = _T_1429 ^ _T_1433; // @[AesSbox.scala 40:63]
  wire  _T_1453 = matrix_1_1[2] ^ _T_1437; // @[AesSbox.scala 40:63]
  wire  _T_1455 = matrix_1_1[7] ^ matrix_1_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_1457 = matrix_1_1[0] ^ _T_1439; // @[AesSbox.scala 40:63]
  wire  _T_1459 = matrix_1_1[1] ^ matrix_1_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_1461 = _T_1427 ^ _T_1459; // @[AesSbox.scala 40:63]
  wire  _T_1463 = _T_1431 ^ _T_1453; // @[AesSbox.scala 40:63]
  wire  _T_1465 = _T_1425 ^ _T_1449; // @[AesSbox.scala 40:63]
  wire  _T_1467 = matrix_1_1[7] ^ _T_1431; // @[AesSbox.scala 40:63]
  wire  _T_1469 = _T_1465 ^ _T_1433; // @[AesSbox.scala 40:63]
  wire  _T_1471 = _T_1465 ^ _T_1437; // @[AesSbox.scala 40:63]
  wire  _T_1473 = _T_1437 ^ _T_1461; // @[AesSbox.scala 40:63]
  wire  _T_1475 = _T_1455 ^ _T_1451; // @[AesSbox.scala 40:63]
  wire  _T_1477 = _T_1467 ^ _T_1457; // @[AesSbox.scala 40:63]
  wire  _T_1479 = _T_1461 & _T_1433; // @[AesSbox.scala 41:63]
  wire  _T_1481 = _T_1463 & _T_1445; // @[AesSbox.scala 41:63]
  wire  _T_1483 = _T_1447 ^ _T_1479; // @[AesSbox.scala 40:63]
  wire  _T_1485 = _T_1443 & matrix_1_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_1487 = _T_1485 ^ _T_1479; // @[AesSbox.scala 40:63]
  wire  _T_1489 = _T_1437 & _T_1465; // @[AesSbox.scala 41:63]
  wire  _T_1491 = _T_1441 & _T_1431; // @[AesSbox.scala 41:63]
  wire  _T_1493 = _T_1471 ^ _T_1489; // @[AesSbox.scala 40:63]
  wire  _T_1495 = _T_1467 & _T_1457; // @[AesSbox.scala 41:63]
  wire  _T_1497 = _T_1495 ^ _T_1489; // @[AesSbox.scala 40:63]
  wire  _T_1499 = _T_1427 & _T_1439; // @[AesSbox.scala 41:63]
  wire  _T_1501 = _T_1473 & _T_1469; // @[AesSbox.scala 41:63]
  wire  _T_1503 = _T_1501 ^ _T_1499; // @[AesSbox.scala 40:63]
  wire  _T_1505 = _T_1455 & _T_1451; // @[AesSbox.scala 41:63]
  wire  _T_1507 = _T_1505 ^ _T_1499; // @[AesSbox.scala 40:63]
  wire  _T_1509 = _T_1483 ^ _T_1481; // @[AesSbox.scala 40:63]
  wire  _T_1511 = _T_1487 ^ _T_1475; // @[AesSbox.scala 40:63]
  wire  _T_1513 = _T_1493 ^ _T_1491; // @[AesSbox.scala 40:63]
  wire  _T_1515 = _T_1497 ^ _T_1507; // @[AesSbox.scala 40:63]
  wire  _T_1517 = _T_1509 ^ _T_1503; // @[AesSbox.scala 40:63]
  wire  _T_1519 = _T_1511 ^ _T_1507; // @[AesSbox.scala 40:63]
  wire  _T_1521 = _T_1513 ^ _T_1503; // @[AesSbox.scala 40:63]
  wire  _T_1523 = _T_1515 ^ _T_1477; // @[AesSbox.scala 40:63]
  wire  _T_1525 = _T_1521 ^ _T_1523; // @[AesSbox.scala 40:63]
  wire  _T_1527 = _T_1521 & _T_1517; // @[AesSbox.scala 41:63]
  wire  _T_1529 = _T_1519 ^ _T_1527; // @[AesSbox.scala 40:63]
  wire  _T_1531 = _T_1517 ^ _T_1519; // @[AesSbox.scala 40:63]
  wire  _T_1533 = _T_1523 ^ _T_1527; // @[AesSbox.scala 40:63]
  wire  _T_1535 = _T_1533 & _T_1531; // @[AesSbox.scala 41:63]
  wire  _T_1537 = _T_1529 & _T_1525; // @[AesSbox.scala 41:63]
  wire  _T_1539 = _T_1517 & _T_1523; // @[AesSbox.scala 41:63]
  wire  _T_1541 = _T_1531 & _T_1539; // @[AesSbox.scala 41:63]
  wire  _T_1543 = _T_1531 ^ _T_1527; // @[AesSbox.scala 40:63]
  wire  _T_1545 = _T_1519 & _T_1521; // @[AesSbox.scala 41:63]
  wire  _T_1547 = _T_1525 & _T_1545; // @[AesSbox.scala 41:63]
  wire  _T_1549 = _T_1525 ^ _T_1527; // @[AesSbox.scala 40:63]
  wire  _T_1551 = _T_1519 ^ _T_1535; // @[AesSbox.scala 40:63]
  wire  _T_1553 = _T_1541 ^ _T_1543; // @[AesSbox.scala 40:63]
  wire  _T_1555 = _T_1523 ^ _T_1537; // @[AesSbox.scala 40:63]
  wire  _T_1557 = _T_1547 ^ _T_1549; // @[AesSbox.scala 40:63]
  wire  _T_1559 = _T_1553 ^ _T_1557; // @[AesSbox.scala 40:63]
  wire  _T_1561 = _T_1551 ^ _T_1555; // @[AesSbox.scala 40:63]
  wire  _T_1563 = _T_1551 ^ _T_1553; // @[AesSbox.scala 40:63]
  wire  _T_1565 = _T_1555 ^ _T_1557; // @[AesSbox.scala 40:63]
  wire  _T_1567 = _T_1561 ^ _T_1559; // @[AesSbox.scala 40:63]
  wire  _T_1569 = _T_1565 & _T_1433; // @[AesSbox.scala 41:63]
  wire  _T_1571 = _T_1557 & _T_1445; // @[AesSbox.scala 41:63]
  wire  _T_1573 = _T_1555 & matrix_1_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_1575 = _T_1563 & _T_1465; // @[AesSbox.scala 41:63]
  wire  _T_1577 = _T_1553 & _T_1431; // @[AesSbox.scala 41:63]
  wire  _T_1579 = _T_1551 & _T_1457; // @[AesSbox.scala 41:63]
  wire  _T_1581 = _T_1561 & _T_1439; // @[AesSbox.scala 41:63]
  wire  _T_1583 = _T_1567 & _T_1469; // @[AesSbox.scala 41:63]
  wire  _T_1585 = _T_1559 & _T_1451; // @[AesSbox.scala 41:63]
  wire  _T_1587 = _T_1565 & _T_1461; // @[AesSbox.scala 41:63]
  wire  _T_1589 = _T_1557 & _T_1463; // @[AesSbox.scala 41:63]
  wire  _T_1591 = _T_1555 & _T_1443; // @[AesSbox.scala 41:63]
  wire  _T_1593 = _T_1563 & _T_1437; // @[AesSbox.scala 41:63]
  wire  _T_1595 = _T_1553 & _T_1441; // @[AesSbox.scala 41:63]
  wire  _T_1597 = _T_1551 & _T_1467; // @[AesSbox.scala 41:63]
  wire  _T_1599 = _T_1561 & _T_1427; // @[AesSbox.scala 41:63]
  wire  _T_1601 = _T_1567 & _T_1473; // @[AesSbox.scala 41:63]
  wire  _T_1603 = _T_1559 & _T_1455; // @[AesSbox.scala 41:63]
  wire  _T_1605 = _T_1599 ^ _T_1601; // @[AesSbox.scala 40:63]
  wire  _T_1607 = _T_1577 ^ _T_1589; // @[AesSbox.scala 40:63]
  wire  _T_1609 = _T_1583 ^ _T_1605; // @[AesSbox.scala 40:63]
  wire  _T_1611 = _T_1587 ^ _T_1607; // @[AesSbox.scala 40:63]
  wire  _T_1613 = _T_1573 ^ _T_1593; // @[AesSbox.scala 40:63]
  wire  _T_1615 = _T_1569 ^ _T_1575; // @[AesSbox.scala 40:63]
  wire  _T_1617 = _T_1605 ^ _T_1615; // @[AesSbox.scala 40:63]
  wire  _T_1619 = _T_1571 ^ _T_1611; // @[AesSbox.scala 40:63]
  wire  _T_1621 = _T_1569 ^ _T_1581; // @[AesSbox.scala 40:63]
  wire  _T_1623 = _T_1579 ^ _T_1595; // @[AesSbox.scala 40:63]
  wire  _T_1625 = _T_1585 ^ _T_1597; // @[AesSbox.scala 40:63]
  wire  _T_1627 = _T_1573 ^ _T_1619; // @[AesSbox.scala 40:63]
  wire  _T_1629 = _T_1613 ^ _T_1625; // @[AesSbox.scala 40:63]
  wire  _T_1631 = _T_1591 ^ _T_1607; // @[AesSbox.scala 40:63]
  wire  _T_1633 = _T_1575 ^ _T_1581; // @[AesSbox.scala 40:63]
  wire  _T_1635 = _T_1611 ^ _T_1633; // @[AesSbox.scala 40:63]
  wire  _T_1637 = _T_1603 ^ _T_1629; // @[AesSbox.scala 40:63]
  wire  _T_1639 = _T_1599 ^ _T_1621; // @[AesSbox.scala 40:63]
  wire  _T_1641 = _T_1613 ^ _T_1623; // @[AesSbox.scala 40:63]
  wire  _T_1642 = _T_1609 ^ _T_1635; // @[AesSbox.scala 40:63]
  wire  _T_1643 = _T_1637 ^ _T_1639; // @[AesSbox.scala 42:65]
  wire  _T_1644 = ~_T_1643; // @[AesSbox.scala 42:51]
  wire  _T_1646 = _T_1579 ^ _T_1605; // @[AesSbox.scala 40:63]
  wire  _T_1647 = _T_1617 ^ _T_1619; // @[AesSbox.scala 40:63]
  wire  _T_1648 = _T_1627 ^ _T_1646; // @[AesSbox.scala 40:63]
  wire  _T_1650 = _T_1577 ^ _T_1593; // @[AesSbox.scala 40:63]
  wire  _T_1652 = _T_1615 ^ _T_1631; // @[AesSbox.scala 40:63]
  wire  _T_1653 = _T_1617 ^ _T_1641; // @[AesSbox.scala 42:65]
  wire  _T_1654 = ~_T_1653; // @[AesSbox.scala 42:51]
  wire  _T_1656 = _T_1585 ^ _T_1623; // @[AesSbox.scala 40:63]
  wire  _T_1658 = _T_1650 ^ _T_1656; // @[AesSbox.scala 40:63]
  wire  _T_1660 = _T_1577 ^ _T_1621; // @[AesSbox.scala 40:63]
  wire  _T_1661 = _T_1609 ^ _T_1658; // @[AesSbox.scala 42:65]
  wire  _T_1662 = ~_T_1661; // @[AesSbox.scala 42:51]
  wire  _T_1664 = _T_1629 ^ _T_1652; // @[AesSbox.scala 40:63]
  wire  _T_1665 = _T_1609 ^ _T_1664; // @[AesSbox.scala 40:63]
  wire  _T_1667 = _T_1619 ^ _T_1660; // @[AesSbox.scala 40:63]
  wire  _T_1668 = _T_1609 ^ _T_1667; // @[AesSbox.scala 42:65]
  wire  _T_1669 = ~_T_1668; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_0_1 = {_T_1642,_T_1669,_T_1644,_T_1647,_T_1648,_T_1665,_T_1662,_T_1654}; // @[Cat.scala 29:58]
  wire  _T_1694 = matrix_1_2[1] ^ matrix_1_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_1696 = matrix_1_2[4] ^ matrix_1_2[7]; // @[AesSbox.scala 40:63]
  wire  _T_1698 = matrix_1_2[6] ^ matrix_1_2[5]; // @[AesSbox.scala 40:63]
  wire  _T_1700 = matrix_1_2[0] ^ _T_1698; // @[AesSbox.scala 40:63]
  wire  _T_1702 = _T_1694 ^ _T_1696; // @[AesSbox.scala 40:63]
  wire  _T_1704 = matrix_1_2[6] ^ matrix_1_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_1706 = matrix_1_2[7] ^ matrix_1_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_1708 = _T_1694 ^ _T_1704; // @[AesSbox.scala 40:63]
  wire  _T_1710 = matrix_1_2[1] ^ _T_1700; // @[AesSbox.scala 40:63]
  wire  _T_1712 = matrix_1_2[4] ^ _T_1700; // @[AesSbox.scala 40:63]
  wire  _T_1714 = matrix_1_2[0] ^ _T_1702; // @[AesSbox.scala 40:63]
  wire  _T_1716 = _T_1702 ^ _T_1704; // @[AesSbox.scala 40:63]
  wire  _T_1718 = matrix_1_2[5] ^ matrix_1_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_1720 = _T_1698 ^ _T_1702; // @[AesSbox.scala 40:63]
  wire  _T_1722 = matrix_1_2[2] ^ _T_1706; // @[AesSbox.scala 40:63]
  wire  _T_1724 = matrix_1_2[7] ^ matrix_1_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_1726 = matrix_1_2[0] ^ _T_1708; // @[AesSbox.scala 40:63]
  wire  _T_1728 = matrix_1_2[1] ^ matrix_1_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_1730 = _T_1696 ^ _T_1728; // @[AesSbox.scala 40:63]
  wire  _T_1732 = _T_1700 ^ _T_1722; // @[AesSbox.scala 40:63]
  wire  _T_1734 = _T_1694 ^ _T_1718; // @[AesSbox.scala 40:63]
  wire  _T_1736 = matrix_1_2[7] ^ _T_1700; // @[AesSbox.scala 40:63]
  wire  _T_1738 = _T_1734 ^ _T_1702; // @[AesSbox.scala 40:63]
  wire  _T_1740 = _T_1734 ^ _T_1706; // @[AesSbox.scala 40:63]
  wire  _T_1742 = _T_1706 ^ _T_1730; // @[AesSbox.scala 40:63]
  wire  _T_1744 = _T_1724 ^ _T_1720; // @[AesSbox.scala 40:63]
  wire  _T_1746 = _T_1736 ^ _T_1726; // @[AesSbox.scala 40:63]
  wire  _T_1748 = _T_1730 & _T_1702; // @[AesSbox.scala 41:63]
  wire  _T_1750 = _T_1732 & _T_1714; // @[AesSbox.scala 41:63]
  wire  _T_1752 = _T_1716 ^ _T_1748; // @[AesSbox.scala 40:63]
  wire  _T_1754 = _T_1712 & matrix_1_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_1756 = _T_1754 ^ _T_1748; // @[AesSbox.scala 40:63]
  wire  _T_1758 = _T_1706 & _T_1734; // @[AesSbox.scala 41:63]
  wire  _T_1760 = _T_1710 & _T_1700; // @[AesSbox.scala 41:63]
  wire  _T_1762 = _T_1740 ^ _T_1758; // @[AesSbox.scala 40:63]
  wire  _T_1764 = _T_1736 & _T_1726; // @[AesSbox.scala 41:63]
  wire  _T_1766 = _T_1764 ^ _T_1758; // @[AesSbox.scala 40:63]
  wire  _T_1768 = _T_1696 & _T_1708; // @[AesSbox.scala 41:63]
  wire  _T_1770 = _T_1742 & _T_1738; // @[AesSbox.scala 41:63]
  wire  _T_1772 = _T_1770 ^ _T_1768; // @[AesSbox.scala 40:63]
  wire  _T_1774 = _T_1724 & _T_1720; // @[AesSbox.scala 41:63]
  wire  _T_1776 = _T_1774 ^ _T_1768; // @[AesSbox.scala 40:63]
  wire  _T_1778 = _T_1752 ^ _T_1750; // @[AesSbox.scala 40:63]
  wire  _T_1780 = _T_1756 ^ _T_1744; // @[AesSbox.scala 40:63]
  wire  _T_1782 = _T_1762 ^ _T_1760; // @[AesSbox.scala 40:63]
  wire  _T_1784 = _T_1766 ^ _T_1776; // @[AesSbox.scala 40:63]
  wire  _T_1786 = _T_1778 ^ _T_1772; // @[AesSbox.scala 40:63]
  wire  _T_1788 = _T_1780 ^ _T_1776; // @[AesSbox.scala 40:63]
  wire  _T_1790 = _T_1782 ^ _T_1772; // @[AesSbox.scala 40:63]
  wire  _T_1792 = _T_1784 ^ _T_1746; // @[AesSbox.scala 40:63]
  wire  _T_1794 = _T_1790 ^ _T_1792; // @[AesSbox.scala 40:63]
  wire  _T_1796 = _T_1790 & _T_1786; // @[AesSbox.scala 41:63]
  wire  _T_1798 = _T_1788 ^ _T_1796; // @[AesSbox.scala 40:63]
  wire  _T_1800 = _T_1786 ^ _T_1788; // @[AesSbox.scala 40:63]
  wire  _T_1802 = _T_1792 ^ _T_1796; // @[AesSbox.scala 40:63]
  wire  _T_1804 = _T_1802 & _T_1800; // @[AesSbox.scala 41:63]
  wire  _T_1806 = _T_1798 & _T_1794; // @[AesSbox.scala 41:63]
  wire  _T_1808 = _T_1786 & _T_1792; // @[AesSbox.scala 41:63]
  wire  _T_1810 = _T_1800 & _T_1808; // @[AesSbox.scala 41:63]
  wire  _T_1812 = _T_1800 ^ _T_1796; // @[AesSbox.scala 40:63]
  wire  _T_1814 = _T_1788 & _T_1790; // @[AesSbox.scala 41:63]
  wire  _T_1816 = _T_1794 & _T_1814; // @[AesSbox.scala 41:63]
  wire  _T_1818 = _T_1794 ^ _T_1796; // @[AesSbox.scala 40:63]
  wire  _T_1820 = _T_1788 ^ _T_1804; // @[AesSbox.scala 40:63]
  wire  _T_1822 = _T_1810 ^ _T_1812; // @[AesSbox.scala 40:63]
  wire  _T_1824 = _T_1792 ^ _T_1806; // @[AesSbox.scala 40:63]
  wire  _T_1826 = _T_1816 ^ _T_1818; // @[AesSbox.scala 40:63]
  wire  _T_1828 = _T_1822 ^ _T_1826; // @[AesSbox.scala 40:63]
  wire  _T_1830 = _T_1820 ^ _T_1824; // @[AesSbox.scala 40:63]
  wire  _T_1832 = _T_1820 ^ _T_1822; // @[AesSbox.scala 40:63]
  wire  _T_1834 = _T_1824 ^ _T_1826; // @[AesSbox.scala 40:63]
  wire  _T_1836 = _T_1830 ^ _T_1828; // @[AesSbox.scala 40:63]
  wire  _T_1838 = _T_1834 & _T_1702; // @[AesSbox.scala 41:63]
  wire  _T_1840 = _T_1826 & _T_1714; // @[AesSbox.scala 41:63]
  wire  _T_1842 = _T_1824 & matrix_1_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_1844 = _T_1832 & _T_1734; // @[AesSbox.scala 41:63]
  wire  _T_1846 = _T_1822 & _T_1700; // @[AesSbox.scala 41:63]
  wire  _T_1848 = _T_1820 & _T_1726; // @[AesSbox.scala 41:63]
  wire  _T_1850 = _T_1830 & _T_1708; // @[AesSbox.scala 41:63]
  wire  _T_1852 = _T_1836 & _T_1738; // @[AesSbox.scala 41:63]
  wire  _T_1854 = _T_1828 & _T_1720; // @[AesSbox.scala 41:63]
  wire  _T_1856 = _T_1834 & _T_1730; // @[AesSbox.scala 41:63]
  wire  _T_1858 = _T_1826 & _T_1732; // @[AesSbox.scala 41:63]
  wire  _T_1860 = _T_1824 & _T_1712; // @[AesSbox.scala 41:63]
  wire  _T_1862 = _T_1832 & _T_1706; // @[AesSbox.scala 41:63]
  wire  _T_1864 = _T_1822 & _T_1710; // @[AesSbox.scala 41:63]
  wire  _T_1866 = _T_1820 & _T_1736; // @[AesSbox.scala 41:63]
  wire  _T_1868 = _T_1830 & _T_1696; // @[AesSbox.scala 41:63]
  wire  _T_1870 = _T_1836 & _T_1742; // @[AesSbox.scala 41:63]
  wire  _T_1872 = _T_1828 & _T_1724; // @[AesSbox.scala 41:63]
  wire  _T_1874 = _T_1868 ^ _T_1870; // @[AesSbox.scala 40:63]
  wire  _T_1876 = _T_1846 ^ _T_1858; // @[AesSbox.scala 40:63]
  wire  _T_1878 = _T_1852 ^ _T_1874; // @[AesSbox.scala 40:63]
  wire  _T_1880 = _T_1856 ^ _T_1876; // @[AesSbox.scala 40:63]
  wire  _T_1882 = _T_1842 ^ _T_1862; // @[AesSbox.scala 40:63]
  wire  _T_1884 = _T_1838 ^ _T_1844; // @[AesSbox.scala 40:63]
  wire  _T_1886 = _T_1874 ^ _T_1884; // @[AesSbox.scala 40:63]
  wire  _T_1888 = _T_1840 ^ _T_1880; // @[AesSbox.scala 40:63]
  wire  _T_1890 = _T_1838 ^ _T_1850; // @[AesSbox.scala 40:63]
  wire  _T_1892 = _T_1848 ^ _T_1864; // @[AesSbox.scala 40:63]
  wire  _T_1894 = _T_1854 ^ _T_1866; // @[AesSbox.scala 40:63]
  wire  _T_1896 = _T_1842 ^ _T_1888; // @[AesSbox.scala 40:63]
  wire  _T_1898 = _T_1882 ^ _T_1894; // @[AesSbox.scala 40:63]
  wire  _T_1900 = _T_1860 ^ _T_1876; // @[AesSbox.scala 40:63]
  wire  _T_1902 = _T_1844 ^ _T_1850; // @[AesSbox.scala 40:63]
  wire  _T_1904 = _T_1880 ^ _T_1902; // @[AesSbox.scala 40:63]
  wire  _T_1906 = _T_1872 ^ _T_1898; // @[AesSbox.scala 40:63]
  wire  _T_1908 = _T_1868 ^ _T_1890; // @[AesSbox.scala 40:63]
  wire  _T_1910 = _T_1882 ^ _T_1892; // @[AesSbox.scala 40:63]
  wire  _T_1911 = _T_1878 ^ _T_1904; // @[AesSbox.scala 40:63]
  wire  _T_1912 = _T_1906 ^ _T_1908; // @[AesSbox.scala 42:65]
  wire  _T_1913 = ~_T_1912; // @[AesSbox.scala 42:51]
  wire  _T_1915 = _T_1848 ^ _T_1874; // @[AesSbox.scala 40:63]
  wire  _T_1916 = _T_1886 ^ _T_1888; // @[AesSbox.scala 40:63]
  wire  _T_1917 = _T_1896 ^ _T_1915; // @[AesSbox.scala 40:63]
  wire  _T_1919 = _T_1846 ^ _T_1862; // @[AesSbox.scala 40:63]
  wire  _T_1921 = _T_1884 ^ _T_1900; // @[AesSbox.scala 40:63]
  wire  _T_1922 = _T_1886 ^ _T_1910; // @[AesSbox.scala 42:65]
  wire  _T_1923 = ~_T_1922; // @[AesSbox.scala 42:51]
  wire  _T_1925 = _T_1854 ^ _T_1892; // @[AesSbox.scala 40:63]
  wire  _T_1927 = _T_1919 ^ _T_1925; // @[AesSbox.scala 40:63]
  wire  _T_1929 = _T_1846 ^ _T_1890; // @[AesSbox.scala 40:63]
  wire  _T_1930 = _T_1878 ^ _T_1927; // @[AesSbox.scala 42:65]
  wire  _T_1931 = ~_T_1930; // @[AesSbox.scala 42:51]
  wire  _T_1933 = _T_1898 ^ _T_1921; // @[AesSbox.scala 40:63]
  wire  _T_1934 = _T_1878 ^ _T_1933; // @[AesSbox.scala 40:63]
  wire  _T_1936 = _T_1888 ^ _T_1929; // @[AesSbox.scala 40:63]
  wire  _T_1937 = _T_1878 ^ _T_1936; // @[AesSbox.scala 42:65]
  wire  _T_1938 = ~_T_1937; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_3_2 = {_T_1911,_T_1938,_T_1913,_T_1916,_T_1917,_T_1934,_T_1931,_T_1923}; // @[Cat.scala 29:58]
  wire  _T_1963 = matrix_1_3[1] ^ matrix_1_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_1965 = matrix_1_3[4] ^ matrix_1_3[7]; // @[AesSbox.scala 40:63]
  wire  _T_1967 = matrix_1_3[6] ^ matrix_1_3[5]; // @[AesSbox.scala 40:63]
  wire  _T_1969 = matrix_1_3[0] ^ _T_1967; // @[AesSbox.scala 40:63]
  wire  _T_1971 = _T_1963 ^ _T_1965; // @[AesSbox.scala 40:63]
  wire  _T_1973 = matrix_1_3[6] ^ matrix_1_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_1975 = matrix_1_3[7] ^ matrix_1_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_1977 = _T_1963 ^ _T_1973; // @[AesSbox.scala 40:63]
  wire  _T_1979 = matrix_1_3[1] ^ _T_1969; // @[AesSbox.scala 40:63]
  wire  _T_1981 = matrix_1_3[4] ^ _T_1969; // @[AesSbox.scala 40:63]
  wire  _T_1983 = matrix_1_3[0] ^ _T_1971; // @[AesSbox.scala 40:63]
  wire  _T_1985 = _T_1971 ^ _T_1973; // @[AesSbox.scala 40:63]
  wire  _T_1987 = matrix_1_3[5] ^ matrix_1_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_1989 = _T_1967 ^ _T_1971; // @[AesSbox.scala 40:63]
  wire  _T_1991 = matrix_1_3[2] ^ _T_1975; // @[AesSbox.scala 40:63]
  wire  _T_1993 = matrix_1_3[7] ^ matrix_1_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_1995 = matrix_1_3[0] ^ _T_1977; // @[AesSbox.scala 40:63]
  wire  _T_1997 = matrix_1_3[1] ^ matrix_1_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_1999 = _T_1965 ^ _T_1997; // @[AesSbox.scala 40:63]
  wire  _T_2001 = _T_1969 ^ _T_1991; // @[AesSbox.scala 40:63]
  wire  _T_2003 = _T_1963 ^ _T_1987; // @[AesSbox.scala 40:63]
  wire  _T_2005 = matrix_1_3[7] ^ _T_1969; // @[AesSbox.scala 40:63]
  wire  _T_2007 = _T_2003 ^ _T_1971; // @[AesSbox.scala 40:63]
  wire  _T_2009 = _T_2003 ^ _T_1975; // @[AesSbox.scala 40:63]
  wire  _T_2011 = _T_1975 ^ _T_1999; // @[AesSbox.scala 40:63]
  wire  _T_2013 = _T_1993 ^ _T_1989; // @[AesSbox.scala 40:63]
  wire  _T_2015 = _T_2005 ^ _T_1995; // @[AesSbox.scala 40:63]
  wire  _T_2017 = _T_1999 & _T_1971; // @[AesSbox.scala 41:63]
  wire  _T_2019 = _T_2001 & _T_1983; // @[AesSbox.scala 41:63]
  wire  _T_2021 = _T_1985 ^ _T_2017; // @[AesSbox.scala 40:63]
  wire  _T_2023 = _T_1981 & matrix_1_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_2025 = _T_2023 ^ _T_2017; // @[AesSbox.scala 40:63]
  wire  _T_2027 = _T_1975 & _T_2003; // @[AesSbox.scala 41:63]
  wire  _T_2029 = _T_1979 & _T_1969; // @[AesSbox.scala 41:63]
  wire  _T_2031 = _T_2009 ^ _T_2027; // @[AesSbox.scala 40:63]
  wire  _T_2033 = _T_2005 & _T_1995; // @[AesSbox.scala 41:63]
  wire  _T_2035 = _T_2033 ^ _T_2027; // @[AesSbox.scala 40:63]
  wire  _T_2037 = _T_1965 & _T_1977; // @[AesSbox.scala 41:63]
  wire  _T_2039 = _T_2011 & _T_2007; // @[AesSbox.scala 41:63]
  wire  _T_2041 = _T_2039 ^ _T_2037; // @[AesSbox.scala 40:63]
  wire  _T_2043 = _T_1993 & _T_1989; // @[AesSbox.scala 41:63]
  wire  _T_2045 = _T_2043 ^ _T_2037; // @[AesSbox.scala 40:63]
  wire  _T_2047 = _T_2021 ^ _T_2019; // @[AesSbox.scala 40:63]
  wire  _T_2049 = _T_2025 ^ _T_2013; // @[AesSbox.scala 40:63]
  wire  _T_2051 = _T_2031 ^ _T_2029; // @[AesSbox.scala 40:63]
  wire  _T_2053 = _T_2035 ^ _T_2045; // @[AesSbox.scala 40:63]
  wire  _T_2055 = _T_2047 ^ _T_2041; // @[AesSbox.scala 40:63]
  wire  _T_2057 = _T_2049 ^ _T_2045; // @[AesSbox.scala 40:63]
  wire  _T_2059 = _T_2051 ^ _T_2041; // @[AesSbox.scala 40:63]
  wire  _T_2061 = _T_2053 ^ _T_2015; // @[AesSbox.scala 40:63]
  wire  _T_2063 = _T_2059 ^ _T_2061; // @[AesSbox.scala 40:63]
  wire  _T_2065 = _T_2059 & _T_2055; // @[AesSbox.scala 41:63]
  wire  _T_2067 = _T_2057 ^ _T_2065; // @[AesSbox.scala 40:63]
  wire  _T_2069 = _T_2055 ^ _T_2057; // @[AesSbox.scala 40:63]
  wire  _T_2071 = _T_2061 ^ _T_2065; // @[AesSbox.scala 40:63]
  wire  _T_2073 = _T_2071 & _T_2069; // @[AesSbox.scala 41:63]
  wire  _T_2075 = _T_2067 & _T_2063; // @[AesSbox.scala 41:63]
  wire  _T_2077 = _T_2055 & _T_2061; // @[AesSbox.scala 41:63]
  wire  _T_2079 = _T_2069 & _T_2077; // @[AesSbox.scala 41:63]
  wire  _T_2081 = _T_2069 ^ _T_2065; // @[AesSbox.scala 40:63]
  wire  _T_2083 = _T_2057 & _T_2059; // @[AesSbox.scala 41:63]
  wire  _T_2085 = _T_2063 & _T_2083; // @[AesSbox.scala 41:63]
  wire  _T_2087 = _T_2063 ^ _T_2065; // @[AesSbox.scala 40:63]
  wire  _T_2089 = _T_2057 ^ _T_2073; // @[AesSbox.scala 40:63]
  wire  _T_2091 = _T_2079 ^ _T_2081; // @[AesSbox.scala 40:63]
  wire  _T_2093 = _T_2061 ^ _T_2075; // @[AesSbox.scala 40:63]
  wire  _T_2095 = _T_2085 ^ _T_2087; // @[AesSbox.scala 40:63]
  wire  _T_2097 = _T_2091 ^ _T_2095; // @[AesSbox.scala 40:63]
  wire  _T_2099 = _T_2089 ^ _T_2093; // @[AesSbox.scala 40:63]
  wire  _T_2101 = _T_2089 ^ _T_2091; // @[AesSbox.scala 40:63]
  wire  _T_2103 = _T_2093 ^ _T_2095; // @[AesSbox.scala 40:63]
  wire  _T_2105 = _T_2099 ^ _T_2097; // @[AesSbox.scala 40:63]
  wire  _T_2107 = _T_2103 & _T_1971; // @[AesSbox.scala 41:63]
  wire  _T_2109 = _T_2095 & _T_1983; // @[AesSbox.scala 41:63]
  wire  _T_2111 = _T_2093 & matrix_1_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_2113 = _T_2101 & _T_2003; // @[AesSbox.scala 41:63]
  wire  _T_2115 = _T_2091 & _T_1969; // @[AesSbox.scala 41:63]
  wire  _T_2117 = _T_2089 & _T_1995; // @[AesSbox.scala 41:63]
  wire  _T_2119 = _T_2099 & _T_1977; // @[AesSbox.scala 41:63]
  wire  _T_2121 = _T_2105 & _T_2007; // @[AesSbox.scala 41:63]
  wire  _T_2123 = _T_2097 & _T_1989; // @[AesSbox.scala 41:63]
  wire  _T_2125 = _T_2103 & _T_1999; // @[AesSbox.scala 41:63]
  wire  _T_2127 = _T_2095 & _T_2001; // @[AesSbox.scala 41:63]
  wire  _T_2129 = _T_2093 & _T_1981; // @[AesSbox.scala 41:63]
  wire  _T_2131 = _T_2101 & _T_1975; // @[AesSbox.scala 41:63]
  wire  _T_2133 = _T_2091 & _T_1979; // @[AesSbox.scala 41:63]
  wire  _T_2135 = _T_2089 & _T_2005; // @[AesSbox.scala 41:63]
  wire  _T_2137 = _T_2099 & _T_1965; // @[AesSbox.scala 41:63]
  wire  _T_2139 = _T_2105 & _T_2011; // @[AesSbox.scala 41:63]
  wire  _T_2141 = _T_2097 & _T_1993; // @[AesSbox.scala 41:63]
  wire  _T_2143 = _T_2137 ^ _T_2139; // @[AesSbox.scala 40:63]
  wire  _T_2145 = _T_2115 ^ _T_2127; // @[AesSbox.scala 40:63]
  wire  _T_2147 = _T_2121 ^ _T_2143; // @[AesSbox.scala 40:63]
  wire  _T_2149 = _T_2125 ^ _T_2145; // @[AesSbox.scala 40:63]
  wire  _T_2151 = _T_2111 ^ _T_2131; // @[AesSbox.scala 40:63]
  wire  _T_2153 = _T_2107 ^ _T_2113; // @[AesSbox.scala 40:63]
  wire  _T_2155 = _T_2143 ^ _T_2153; // @[AesSbox.scala 40:63]
  wire  _T_2157 = _T_2109 ^ _T_2149; // @[AesSbox.scala 40:63]
  wire  _T_2159 = _T_2107 ^ _T_2119; // @[AesSbox.scala 40:63]
  wire  _T_2161 = _T_2117 ^ _T_2133; // @[AesSbox.scala 40:63]
  wire  _T_2163 = _T_2123 ^ _T_2135; // @[AesSbox.scala 40:63]
  wire  _T_2165 = _T_2111 ^ _T_2157; // @[AesSbox.scala 40:63]
  wire  _T_2167 = _T_2151 ^ _T_2163; // @[AesSbox.scala 40:63]
  wire  _T_2169 = _T_2129 ^ _T_2145; // @[AesSbox.scala 40:63]
  wire  _T_2171 = _T_2113 ^ _T_2119; // @[AesSbox.scala 40:63]
  wire  _T_2173 = _T_2149 ^ _T_2171; // @[AesSbox.scala 40:63]
  wire  _T_2175 = _T_2141 ^ _T_2167; // @[AesSbox.scala 40:63]
  wire  _T_2177 = _T_2137 ^ _T_2159; // @[AesSbox.scala 40:63]
  wire  _T_2179 = _T_2151 ^ _T_2161; // @[AesSbox.scala 40:63]
  wire  _T_2180 = _T_2147 ^ _T_2173; // @[AesSbox.scala 40:63]
  wire  _T_2181 = _T_2175 ^ _T_2177; // @[AesSbox.scala 42:65]
  wire  _T_2182 = ~_T_2181; // @[AesSbox.scala 42:51]
  wire  _T_2184 = _T_2117 ^ _T_2143; // @[AesSbox.scala 40:63]
  wire  _T_2185 = _T_2155 ^ _T_2157; // @[AesSbox.scala 40:63]
  wire  _T_2186 = _T_2165 ^ _T_2184; // @[AesSbox.scala 40:63]
  wire  _T_2188 = _T_2115 ^ _T_2131; // @[AesSbox.scala 40:63]
  wire  _T_2190 = _T_2153 ^ _T_2169; // @[AesSbox.scala 40:63]
  wire  _T_2191 = _T_2155 ^ _T_2179; // @[AesSbox.scala 42:65]
  wire  _T_2192 = ~_T_2191; // @[AesSbox.scala 42:51]
  wire  _T_2194 = _T_2123 ^ _T_2161; // @[AesSbox.scala 40:63]
  wire  _T_2196 = _T_2188 ^ _T_2194; // @[AesSbox.scala 40:63]
  wire  _T_2198 = _T_2115 ^ _T_2159; // @[AesSbox.scala 40:63]
  wire  _T_2199 = _T_2147 ^ _T_2196; // @[AesSbox.scala 42:65]
  wire  _T_2200 = ~_T_2199; // @[AesSbox.scala 42:51]
  wire  _T_2202 = _T_2167 ^ _T_2190; // @[AesSbox.scala 40:63]
  wire  _T_2203 = _T_2147 ^ _T_2202; // @[AesSbox.scala 40:63]
  wire  _T_2205 = _T_2157 ^ _T_2198; // @[AesSbox.scala 40:63]
  wire  _T_2206 = _T_2147 ^ _T_2205; // @[AesSbox.scala 42:65]
  wire  _T_2207 = ~_T_2206; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_2_3 = {_T_2180,_T_2207,_T_2182,_T_2185,_T_2186,_T_2203,_T_2200,_T_2192}; // @[Cat.scala 29:58]
  wire  _T_2233 = matrix_2_0[1] ^ matrix_2_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_2235 = matrix_2_0[4] ^ matrix_2_0[7]; // @[AesSbox.scala 40:63]
  wire  _T_2237 = matrix_2_0[6] ^ matrix_2_0[5]; // @[AesSbox.scala 40:63]
  wire  _T_2239 = matrix_2_0[0] ^ _T_2237; // @[AesSbox.scala 40:63]
  wire  _T_2241 = _T_2233 ^ _T_2235; // @[AesSbox.scala 40:63]
  wire  _T_2243 = matrix_2_0[6] ^ matrix_2_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_2245 = matrix_2_0[7] ^ matrix_2_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_2247 = _T_2233 ^ _T_2243; // @[AesSbox.scala 40:63]
  wire  _T_2249 = matrix_2_0[1] ^ _T_2239; // @[AesSbox.scala 40:63]
  wire  _T_2251 = matrix_2_0[4] ^ _T_2239; // @[AesSbox.scala 40:63]
  wire  _T_2253 = matrix_2_0[0] ^ _T_2241; // @[AesSbox.scala 40:63]
  wire  _T_2255 = _T_2241 ^ _T_2243; // @[AesSbox.scala 40:63]
  wire  _T_2257 = matrix_2_0[5] ^ matrix_2_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_2259 = _T_2237 ^ _T_2241; // @[AesSbox.scala 40:63]
  wire  _T_2261 = matrix_2_0[2] ^ _T_2245; // @[AesSbox.scala 40:63]
  wire  _T_2263 = matrix_2_0[7] ^ matrix_2_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_2265 = matrix_2_0[0] ^ _T_2247; // @[AesSbox.scala 40:63]
  wire  _T_2267 = matrix_2_0[1] ^ matrix_2_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_2269 = _T_2235 ^ _T_2267; // @[AesSbox.scala 40:63]
  wire  _T_2271 = _T_2239 ^ _T_2261; // @[AesSbox.scala 40:63]
  wire  _T_2273 = _T_2233 ^ _T_2257; // @[AesSbox.scala 40:63]
  wire  _T_2275 = matrix_2_0[7] ^ _T_2239; // @[AesSbox.scala 40:63]
  wire  _T_2277 = _T_2273 ^ _T_2241; // @[AesSbox.scala 40:63]
  wire  _T_2279 = _T_2273 ^ _T_2245; // @[AesSbox.scala 40:63]
  wire  _T_2281 = _T_2245 ^ _T_2269; // @[AesSbox.scala 40:63]
  wire  _T_2283 = _T_2263 ^ _T_2259; // @[AesSbox.scala 40:63]
  wire  _T_2285 = _T_2275 ^ _T_2265; // @[AesSbox.scala 40:63]
  wire  _T_2287 = _T_2269 & _T_2241; // @[AesSbox.scala 41:63]
  wire  _T_2289 = _T_2271 & _T_2253; // @[AesSbox.scala 41:63]
  wire  _T_2291 = _T_2255 ^ _T_2287; // @[AesSbox.scala 40:63]
  wire  _T_2293 = _T_2251 & matrix_2_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_2295 = _T_2293 ^ _T_2287; // @[AesSbox.scala 40:63]
  wire  _T_2297 = _T_2245 & _T_2273; // @[AesSbox.scala 41:63]
  wire  _T_2299 = _T_2249 & _T_2239; // @[AesSbox.scala 41:63]
  wire  _T_2301 = _T_2279 ^ _T_2297; // @[AesSbox.scala 40:63]
  wire  _T_2303 = _T_2275 & _T_2265; // @[AesSbox.scala 41:63]
  wire  _T_2305 = _T_2303 ^ _T_2297; // @[AesSbox.scala 40:63]
  wire  _T_2307 = _T_2235 & _T_2247; // @[AesSbox.scala 41:63]
  wire  _T_2309 = _T_2281 & _T_2277; // @[AesSbox.scala 41:63]
  wire  _T_2311 = _T_2309 ^ _T_2307; // @[AesSbox.scala 40:63]
  wire  _T_2313 = _T_2263 & _T_2259; // @[AesSbox.scala 41:63]
  wire  _T_2315 = _T_2313 ^ _T_2307; // @[AesSbox.scala 40:63]
  wire  _T_2317 = _T_2291 ^ _T_2289; // @[AesSbox.scala 40:63]
  wire  _T_2319 = _T_2295 ^ _T_2283; // @[AesSbox.scala 40:63]
  wire  _T_2321 = _T_2301 ^ _T_2299; // @[AesSbox.scala 40:63]
  wire  _T_2323 = _T_2305 ^ _T_2315; // @[AesSbox.scala 40:63]
  wire  _T_2325 = _T_2317 ^ _T_2311; // @[AesSbox.scala 40:63]
  wire  _T_2327 = _T_2319 ^ _T_2315; // @[AesSbox.scala 40:63]
  wire  _T_2329 = _T_2321 ^ _T_2311; // @[AesSbox.scala 40:63]
  wire  _T_2331 = _T_2323 ^ _T_2285; // @[AesSbox.scala 40:63]
  wire  _T_2333 = _T_2329 ^ _T_2331; // @[AesSbox.scala 40:63]
  wire  _T_2335 = _T_2329 & _T_2325; // @[AesSbox.scala 41:63]
  wire  _T_2337 = _T_2327 ^ _T_2335; // @[AesSbox.scala 40:63]
  wire  _T_2339 = _T_2325 ^ _T_2327; // @[AesSbox.scala 40:63]
  wire  _T_2341 = _T_2331 ^ _T_2335; // @[AesSbox.scala 40:63]
  wire  _T_2343 = _T_2341 & _T_2339; // @[AesSbox.scala 41:63]
  wire  _T_2345 = _T_2337 & _T_2333; // @[AesSbox.scala 41:63]
  wire  _T_2347 = _T_2325 & _T_2331; // @[AesSbox.scala 41:63]
  wire  _T_2349 = _T_2339 & _T_2347; // @[AesSbox.scala 41:63]
  wire  _T_2351 = _T_2339 ^ _T_2335; // @[AesSbox.scala 40:63]
  wire  _T_2353 = _T_2327 & _T_2329; // @[AesSbox.scala 41:63]
  wire  _T_2355 = _T_2333 & _T_2353; // @[AesSbox.scala 41:63]
  wire  _T_2357 = _T_2333 ^ _T_2335; // @[AesSbox.scala 40:63]
  wire  _T_2359 = _T_2327 ^ _T_2343; // @[AesSbox.scala 40:63]
  wire  _T_2361 = _T_2349 ^ _T_2351; // @[AesSbox.scala 40:63]
  wire  _T_2363 = _T_2331 ^ _T_2345; // @[AesSbox.scala 40:63]
  wire  _T_2365 = _T_2355 ^ _T_2357; // @[AesSbox.scala 40:63]
  wire  _T_2367 = _T_2361 ^ _T_2365; // @[AesSbox.scala 40:63]
  wire  _T_2369 = _T_2359 ^ _T_2363; // @[AesSbox.scala 40:63]
  wire  _T_2371 = _T_2359 ^ _T_2361; // @[AesSbox.scala 40:63]
  wire  _T_2373 = _T_2363 ^ _T_2365; // @[AesSbox.scala 40:63]
  wire  _T_2375 = _T_2369 ^ _T_2367; // @[AesSbox.scala 40:63]
  wire  _T_2377 = _T_2373 & _T_2241; // @[AesSbox.scala 41:63]
  wire  _T_2379 = _T_2365 & _T_2253; // @[AesSbox.scala 41:63]
  wire  _T_2381 = _T_2363 & matrix_2_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_2383 = _T_2371 & _T_2273; // @[AesSbox.scala 41:63]
  wire  _T_2385 = _T_2361 & _T_2239; // @[AesSbox.scala 41:63]
  wire  _T_2387 = _T_2359 & _T_2265; // @[AesSbox.scala 41:63]
  wire  _T_2389 = _T_2369 & _T_2247; // @[AesSbox.scala 41:63]
  wire  _T_2391 = _T_2375 & _T_2277; // @[AesSbox.scala 41:63]
  wire  _T_2393 = _T_2367 & _T_2259; // @[AesSbox.scala 41:63]
  wire  _T_2395 = _T_2373 & _T_2269; // @[AesSbox.scala 41:63]
  wire  _T_2397 = _T_2365 & _T_2271; // @[AesSbox.scala 41:63]
  wire  _T_2399 = _T_2363 & _T_2251; // @[AesSbox.scala 41:63]
  wire  _T_2401 = _T_2371 & _T_2245; // @[AesSbox.scala 41:63]
  wire  _T_2403 = _T_2361 & _T_2249; // @[AesSbox.scala 41:63]
  wire  _T_2405 = _T_2359 & _T_2275; // @[AesSbox.scala 41:63]
  wire  _T_2407 = _T_2369 & _T_2235; // @[AesSbox.scala 41:63]
  wire  _T_2409 = _T_2375 & _T_2281; // @[AesSbox.scala 41:63]
  wire  _T_2411 = _T_2367 & _T_2263; // @[AesSbox.scala 41:63]
  wire  _T_2413 = _T_2407 ^ _T_2409; // @[AesSbox.scala 40:63]
  wire  _T_2415 = _T_2385 ^ _T_2397; // @[AesSbox.scala 40:63]
  wire  _T_2417 = _T_2391 ^ _T_2413; // @[AesSbox.scala 40:63]
  wire  _T_2419 = _T_2395 ^ _T_2415; // @[AesSbox.scala 40:63]
  wire  _T_2421 = _T_2381 ^ _T_2401; // @[AesSbox.scala 40:63]
  wire  _T_2423 = _T_2377 ^ _T_2383; // @[AesSbox.scala 40:63]
  wire  _T_2425 = _T_2413 ^ _T_2423; // @[AesSbox.scala 40:63]
  wire  _T_2427 = _T_2379 ^ _T_2419; // @[AesSbox.scala 40:63]
  wire  _T_2429 = _T_2377 ^ _T_2389; // @[AesSbox.scala 40:63]
  wire  _T_2431 = _T_2387 ^ _T_2403; // @[AesSbox.scala 40:63]
  wire  _T_2433 = _T_2393 ^ _T_2405; // @[AesSbox.scala 40:63]
  wire  _T_2435 = _T_2381 ^ _T_2427; // @[AesSbox.scala 40:63]
  wire  _T_2437 = _T_2421 ^ _T_2433; // @[AesSbox.scala 40:63]
  wire  _T_2439 = _T_2399 ^ _T_2415; // @[AesSbox.scala 40:63]
  wire  _T_2441 = _T_2383 ^ _T_2389; // @[AesSbox.scala 40:63]
  wire  _T_2443 = _T_2419 ^ _T_2441; // @[AesSbox.scala 40:63]
  wire  _T_2445 = _T_2411 ^ _T_2437; // @[AesSbox.scala 40:63]
  wire  _T_2447 = _T_2407 ^ _T_2429; // @[AesSbox.scala 40:63]
  wire  _T_2449 = _T_2421 ^ _T_2431; // @[AesSbox.scala 40:63]
  wire  _T_2450 = _T_2417 ^ _T_2443; // @[AesSbox.scala 40:63]
  wire  _T_2451 = _T_2445 ^ _T_2447; // @[AesSbox.scala 42:65]
  wire  _T_2452 = ~_T_2451; // @[AesSbox.scala 42:51]
  wire  _T_2454 = _T_2387 ^ _T_2413; // @[AesSbox.scala 40:63]
  wire  _T_2455 = _T_2425 ^ _T_2427; // @[AesSbox.scala 40:63]
  wire  _T_2456 = _T_2435 ^ _T_2454; // @[AesSbox.scala 40:63]
  wire  _T_2458 = _T_2385 ^ _T_2401; // @[AesSbox.scala 40:63]
  wire  _T_2460 = _T_2423 ^ _T_2439; // @[AesSbox.scala 40:63]
  wire  _T_2461 = _T_2425 ^ _T_2449; // @[AesSbox.scala 42:65]
  wire  _T_2462 = ~_T_2461; // @[AesSbox.scala 42:51]
  wire  _T_2464 = _T_2393 ^ _T_2431; // @[AesSbox.scala 40:63]
  wire  _T_2466 = _T_2458 ^ _T_2464; // @[AesSbox.scala 40:63]
  wire  _T_2468 = _T_2385 ^ _T_2429; // @[AesSbox.scala 40:63]
  wire  _T_2469 = _T_2417 ^ _T_2466; // @[AesSbox.scala 42:65]
  wire  _T_2470 = ~_T_2469; // @[AesSbox.scala 42:51]
  wire  _T_2472 = _T_2437 ^ _T_2460; // @[AesSbox.scala 40:63]
  wire  _T_2473 = _T_2417 ^ _T_2472; // @[AesSbox.scala 40:63]
  wire  _T_2475 = _T_2427 ^ _T_2468; // @[AesSbox.scala 40:63]
  wire  _T_2476 = _T_2417 ^ _T_2475; // @[AesSbox.scala 42:65]
  wire  _T_2477 = ~_T_2476; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_2_0 = {_T_2450,_T_2477,_T_2452,_T_2455,_T_2456,_T_2473,_T_2470,_T_2462}; // @[Cat.scala 29:58]
  wire  _T_2502 = matrix_2_1[1] ^ matrix_2_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_2504 = matrix_2_1[4] ^ matrix_2_1[7]; // @[AesSbox.scala 40:63]
  wire  _T_2506 = matrix_2_1[6] ^ matrix_2_1[5]; // @[AesSbox.scala 40:63]
  wire  _T_2508 = matrix_2_1[0] ^ _T_2506; // @[AesSbox.scala 40:63]
  wire  _T_2510 = _T_2502 ^ _T_2504; // @[AesSbox.scala 40:63]
  wire  _T_2512 = matrix_2_1[6] ^ matrix_2_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_2514 = matrix_2_1[7] ^ matrix_2_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_2516 = _T_2502 ^ _T_2512; // @[AesSbox.scala 40:63]
  wire  _T_2518 = matrix_2_1[1] ^ _T_2508; // @[AesSbox.scala 40:63]
  wire  _T_2520 = matrix_2_1[4] ^ _T_2508; // @[AesSbox.scala 40:63]
  wire  _T_2522 = matrix_2_1[0] ^ _T_2510; // @[AesSbox.scala 40:63]
  wire  _T_2524 = _T_2510 ^ _T_2512; // @[AesSbox.scala 40:63]
  wire  _T_2526 = matrix_2_1[5] ^ matrix_2_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_2528 = _T_2506 ^ _T_2510; // @[AesSbox.scala 40:63]
  wire  _T_2530 = matrix_2_1[2] ^ _T_2514; // @[AesSbox.scala 40:63]
  wire  _T_2532 = matrix_2_1[7] ^ matrix_2_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_2534 = matrix_2_1[0] ^ _T_2516; // @[AesSbox.scala 40:63]
  wire  _T_2536 = matrix_2_1[1] ^ matrix_2_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_2538 = _T_2504 ^ _T_2536; // @[AesSbox.scala 40:63]
  wire  _T_2540 = _T_2508 ^ _T_2530; // @[AesSbox.scala 40:63]
  wire  _T_2542 = _T_2502 ^ _T_2526; // @[AesSbox.scala 40:63]
  wire  _T_2544 = matrix_2_1[7] ^ _T_2508; // @[AesSbox.scala 40:63]
  wire  _T_2546 = _T_2542 ^ _T_2510; // @[AesSbox.scala 40:63]
  wire  _T_2548 = _T_2542 ^ _T_2514; // @[AesSbox.scala 40:63]
  wire  _T_2550 = _T_2514 ^ _T_2538; // @[AesSbox.scala 40:63]
  wire  _T_2552 = _T_2532 ^ _T_2528; // @[AesSbox.scala 40:63]
  wire  _T_2554 = _T_2544 ^ _T_2534; // @[AesSbox.scala 40:63]
  wire  _T_2556 = _T_2538 & _T_2510; // @[AesSbox.scala 41:63]
  wire  _T_2558 = _T_2540 & _T_2522; // @[AesSbox.scala 41:63]
  wire  _T_2560 = _T_2524 ^ _T_2556; // @[AesSbox.scala 40:63]
  wire  _T_2562 = _T_2520 & matrix_2_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_2564 = _T_2562 ^ _T_2556; // @[AesSbox.scala 40:63]
  wire  _T_2566 = _T_2514 & _T_2542; // @[AesSbox.scala 41:63]
  wire  _T_2568 = _T_2518 & _T_2508; // @[AesSbox.scala 41:63]
  wire  _T_2570 = _T_2548 ^ _T_2566; // @[AesSbox.scala 40:63]
  wire  _T_2572 = _T_2544 & _T_2534; // @[AesSbox.scala 41:63]
  wire  _T_2574 = _T_2572 ^ _T_2566; // @[AesSbox.scala 40:63]
  wire  _T_2576 = _T_2504 & _T_2516; // @[AesSbox.scala 41:63]
  wire  _T_2578 = _T_2550 & _T_2546; // @[AesSbox.scala 41:63]
  wire  _T_2580 = _T_2578 ^ _T_2576; // @[AesSbox.scala 40:63]
  wire  _T_2582 = _T_2532 & _T_2528; // @[AesSbox.scala 41:63]
  wire  _T_2584 = _T_2582 ^ _T_2576; // @[AesSbox.scala 40:63]
  wire  _T_2586 = _T_2560 ^ _T_2558; // @[AesSbox.scala 40:63]
  wire  _T_2588 = _T_2564 ^ _T_2552; // @[AesSbox.scala 40:63]
  wire  _T_2590 = _T_2570 ^ _T_2568; // @[AesSbox.scala 40:63]
  wire  _T_2592 = _T_2574 ^ _T_2584; // @[AesSbox.scala 40:63]
  wire  _T_2594 = _T_2586 ^ _T_2580; // @[AesSbox.scala 40:63]
  wire  _T_2596 = _T_2588 ^ _T_2584; // @[AesSbox.scala 40:63]
  wire  _T_2598 = _T_2590 ^ _T_2580; // @[AesSbox.scala 40:63]
  wire  _T_2600 = _T_2592 ^ _T_2554; // @[AesSbox.scala 40:63]
  wire  _T_2602 = _T_2598 ^ _T_2600; // @[AesSbox.scala 40:63]
  wire  _T_2604 = _T_2598 & _T_2594; // @[AesSbox.scala 41:63]
  wire  _T_2606 = _T_2596 ^ _T_2604; // @[AesSbox.scala 40:63]
  wire  _T_2608 = _T_2594 ^ _T_2596; // @[AesSbox.scala 40:63]
  wire  _T_2610 = _T_2600 ^ _T_2604; // @[AesSbox.scala 40:63]
  wire  _T_2612 = _T_2610 & _T_2608; // @[AesSbox.scala 41:63]
  wire  _T_2614 = _T_2606 & _T_2602; // @[AesSbox.scala 41:63]
  wire  _T_2616 = _T_2594 & _T_2600; // @[AesSbox.scala 41:63]
  wire  _T_2618 = _T_2608 & _T_2616; // @[AesSbox.scala 41:63]
  wire  _T_2620 = _T_2608 ^ _T_2604; // @[AesSbox.scala 40:63]
  wire  _T_2622 = _T_2596 & _T_2598; // @[AesSbox.scala 41:63]
  wire  _T_2624 = _T_2602 & _T_2622; // @[AesSbox.scala 41:63]
  wire  _T_2626 = _T_2602 ^ _T_2604; // @[AesSbox.scala 40:63]
  wire  _T_2628 = _T_2596 ^ _T_2612; // @[AesSbox.scala 40:63]
  wire  _T_2630 = _T_2618 ^ _T_2620; // @[AesSbox.scala 40:63]
  wire  _T_2632 = _T_2600 ^ _T_2614; // @[AesSbox.scala 40:63]
  wire  _T_2634 = _T_2624 ^ _T_2626; // @[AesSbox.scala 40:63]
  wire  _T_2636 = _T_2630 ^ _T_2634; // @[AesSbox.scala 40:63]
  wire  _T_2638 = _T_2628 ^ _T_2632; // @[AesSbox.scala 40:63]
  wire  _T_2640 = _T_2628 ^ _T_2630; // @[AesSbox.scala 40:63]
  wire  _T_2642 = _T_2632 ^ _T_2634; // @[AesSbox.scala 40:63]
  wire  _T_2644 = _T_2638 ^ _T_2636; // @[AesSbox.scala 40:63]
  wire  _T_2646 = _T_2642 & _T_2510; // @[AesSbox.scala 41:63]
  wire  _T_2648 = _T_2634 & _T_2522; // @[AesSbox.scala 41:63]
  wire  _T_2650 = _T_2632 & matrix_2_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_2652 = _T_2640 & _T_2542; // @[AesSbox.scala 41:63]
  wire  _T_2654 = _T_2630 & _T_2508; // @[AesSbox.scala 41:63]
  wire  _T_2656 = _T_2628 & _T_2534; // @[AesSbox.scala 41:63]
  wire  _T_2658 = _T_2638 & _T_2516; // @[AesSbox.scala 41:63]
  wire  _T_2660 = _T_2644 & _T_2546; // @[AesSbox.scala 41:63]
  wire  _T_2662 = _T_2636 & _T_2528; // @[AesSbox.scala 41:63]
  wire  _T_2664 = _T_2642 & _T_2538; // @[AesSbox.scala 41:63]
  wire  _T_2666 = _T_2634 & _T_2540; // @[AesSbox.scala 41:63]
  wire  _T_2668 = _T_2632 & _T_2520; // @[AesSbox.scala 41:63]
  wire  _T_2670 = _T_2640 & _T_2514; // @[AesSbox.scala 41:63]
  wire  _T_2672 = _T_2630 & _T_2518; // @[AesSbox.scala 41:63]
  wire  _T_2674 = _T_2628 & _T_2544; // @[AesSbox.scala 41:63]
  wire  _T_2676 = _T_2638 & _T_2504; // @[AesSbox.scala 41:63]
  wire  _T_2678 = _T_2644 & _T_2550; // @[AesSbox.scala 41:63]
  wire  _T_2680 = _T_2636 & _T_2532; // @[AesSbox.scala 41:63]
  wire  _T_2682 = _T_2676 ^ _T_2678; // @[AesSbox.scala 40:63]
  wire  _T_2684 = _T_2654 ^ _T_2666; // @[AesSbox.scala 40:63]
  wire  _T_2686 = _T_2660 ^ _T_2682; // @[AesSbox.scala 40:63]
  wire  _T_2688 = _T_2664 ^ _T_2684; // @[AesSbox.scala 40:63]
  wire  _T_2690 = _T_2650 ^ _T_2670; // @[AesSbox.scala 40:63]
  wire  _T_2692 = _T_2646 ^ _T_2652; // @[AesSbox.scala 40:63]
  wire  _T_2694 = _T_2682 ^ _T_2692; // @[AesSbox.scala 40:63]
  wire  _T_2696 = _T_2648 ^ _T_2688; // @[AesSbox.scala 40:63]
  wire  _T_2698 = _T_2646 ^ _T_2658; // @[AesSbox.scala 40:63]
  wire  _T_2700 = _T_2656 ^ _T_2672; // @[AesSbox.scala 40:63]
  wire  _T_2702 = _T_2662 ^ _T_2674; // @[AesSbox.scala 40:63]
  wire  _T_2704 = _T_2650 ^ _T_2696; // @[AesSbox.scala 40:63]
  wire  _T_2706 = _T_2690 ^ _T_2702; // @[AesSbox.scala 40:63]
  wire  _T_2708 = _T_2668 ^ _T_2684; // @[AesSbox.scala 40:63]
  wire  _T_2710 = _T_2652 ^ _T_2658; // @[AesSbox.scala 40:63]
  wire  _T_2712 = _T_2688 ^ _T_2710; // @[AesSbox.scala 40:63]
  wire  _T_2714 = _T_2680 ^ _T_2706; // @[AesSbox.scala 40:63]
  wire  _T_2716 = _T_2676 ^ _T_2698; // @[AesSbox.scala 40:63]
  wire  _T_2718 = _T_2690 ^ _T_2700; // @[AesSbox.scala 40:63]
  wire  _T_2719 = _T_2686 ^ _T_2712; // @[AesSbox.scala 40:63]
  wire  _T_2720 = _T_2714 ^ _T_2716; // @[AesSbox.scala 42:65]
  wire  _T_2721 = ~_T_2720; // @[AesSbox.scala 42:51]
  wire  _T_2723 = _T_2656 ^ _T_2682; // @[AesSbox.scala 40:63]
  wire  _T_2724 = _T_2694 ^ _T_2696; // @[AesSbox.scala 40:63]
  wire  _T_2725 = _T_2704 ^ _T_2723; // @[AesSbox.scala 40:63]
  wire  _T_2727 = _T_2654 ^ _T_2670; // @[AesSbox.scala 40:63]
  wire  _T_2729 = _T_2692 ^ _T_2708; // @[AesSbox.scala 40:63]
  wire  _T_2730 = _T_2694 ^ _T_2718; // @[AesSbox.scala 42:65]
  wire  _T_2731 = ~_T_2730; // @[AesSbox.scala 42:51]
  wire  _T_2733 = _T_2662 ^ _T_2700; // @[AesSbox.scala 40:63]
  wire  _T_2735 = _T_2727 ^ _T_2733; // @[AesSbox.scala 40:63]
  wire  _T_2737 = _T_2654 ^ _T_2698; // @[AesSbox.scala 40:63]
  wire  _T_2738 = _T_2686 ^ _T_2735; // @[AesSbox.scala 42:65]
  wire  _T_2739 = ~_T_2738; // @[AesSbox.scala 42:51]
  wire  _T_2741 = _T_2706 ^ _T_2729; // @[AesSbox.scala 40:63]
  wire  _T_2742 = _T_2686 ^ _T_2741; // @[AesSbox.scala 40:63]
  wire  _T_2744 = _T_2696 ^ _T_2737; // @[AesSbox.scala 40:63]
  wire  _T_2745 = _T_2686 ^ _T_2744; // @[AesSbox.scala 42:65]
  wire  _T_2746 = ~_T_2745; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_1_1 = {_T_2719,_T_2746,_T_2721,_T_2724,_T_2725,_T_2742,_T_2739,_T_2731}; // @[Cat.scala 29:58]
  wire  _T_2771 = matrix_2_2[1] ^ matrix_2_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_2773 = matrix_2_2[4] ^ matrix_2_2[7]; // @[AesSbox.scala 40:63]
  wire  _T_2775 = matrix_2_2[6] ^ matrix_2_2[5]; // @[AesSbox.scala 40:63]
  wire  _T_2777 = matrix_2_2[0] ^ _T_2775; // @[AesSbox.scala 40:63]
  wire  _T_2779 = _T_2771 ^ _T_2773; // @[AesSbox.scala 40:63]
  wire  _T_2781 = matrix_2_2[6] ^ matrix_2_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_2783 = matrix_2_2[7] ^ matrix_2_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_2785 = _T_2771 ^ _T_2781; // @[AesSbox.scala 40:63]
  wire  _T_2787 = matrix_2_2[1] ^ _T_2777; // @[AesSbox.scala 40:63]
  wire  _T_2789 = matrix_2_2[4] ^ _T_2777; // @[AesSbox.scala 40:63]
  wire  _T_2791 = matrix_2_2[0] ^ _T_2779; // @[AesSbox.scala 40:63]
  wire  _T_2793 = _T_2779 ^ _T_2781; // @[AesSbox.scala 40:63]
  wire  _T_2795 = matrix_2_2[5] ^ matrix_2_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_2797 = _T_2775 ^ _T_2779; // @[AesSbox.scala 40:63]
  wire  _T_2799 = matrix_2_2[2] ^ _T_2783; // @[AesSbox.scala 40:63]
  wire  _T_2801 = matrix_2_2[7] ^ matrix_2_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_2803 = matrix_2_2[0] ^ _T_2785; // @[AesSbox.scala 40:63]
  wire  _T_2805 = matrix_2_2[1] ^ matrix_2_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_2807 = _T_2773 ^ _T_2805; // @[AesSbox.scala 40:63]
  wire  _T_2809 = _T_2777 ^ _T_2799; // @[AesSbox.scala 40:63]
  wire  _T_2811 = _T_2771 ^ _T_2795; // @[AesSbox.scala 40:63]
  wire  _T_2813 = matrix_2_2[7] ^ _T_2777; // @[AesSbox.scala 40:63]
  wire  _T_2815 = _T_2811 ^ _T_2779; // @[AesSbox.scala 40:63]
  wire  _T_2817 = _T_2811 ^ _T_2783; // @[AesSbox.scala 40:63]
  wire  _T_2819 = _T_2783 ^ _T_2807; // @[AesSbox.scala 40:63]
  wire  _T_2821 = _T_2801 ^ _T_2797; // @[AesSbox.scala 40:63]
  wire  _T_2823 = _T_2813 ^ _T_2803; // @[AesSbox.scala 40:63]
  wire  _T_2825 = _T_2807 & _T_2779; // @[AesSbox.scala 41:63]
  wire  _T_2827 = _T_2809 & _T_2791; // @[AesSbox.scala 41:63]
  wire  _T_2829 = _T_2793 ^ _T_2825; // @[AesSbox.scala 40:63]
  wire  _T_2831 = _T_2789 & matrix_2_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_2833 = _T_2831 ^ _T_2825; // @[AesSbox.scala 40:63]
  wire  _T_2835 = _T_2783 & _T_2811; // @[AesSbox.scala 41:63]
  wire  _T_2837 = _T_2787 & _T_2777; // @[AesSbox.scala 41:63]
  wire  _T_2839 = _T_2817 ^ _T_2835; // @[AesSbox.scala 40:63]
  wire  _T_2841 = _T_2813 & _T_2803; // @[AesSbox.scala 41:63]
  wire  _T_2843 = _T_2841 ^ _T_2835; // @[AesSbox.scala 40:63]
  wire  _T_2845 = _T_2773 & _T_2785; // @[AesSbox.scala 41:63]
  wire  _T_2847 = _T_2819 & _T_2815; // @[AesSbox.scala 41:63]
  wire  _T_2849 = _T_2847 ^ _T_2845; // @[AesSbox.scala 40:63]
  wire  _T_2851 = _T_2801 & _T_2797; // @[AesSbox.scala 41:63]
  wire  _T_2853 = _T_2851 ^ _T_2845; // @[AesSbox.scala 40:63]
  wire  _T_2855 = _T_2829 ^ _T_2827; // @[AesSbox.scala 40:63]
  wire  _T_2857 = _T_2833 ^ _T_2821; // @[AesSbox.scala 40:63]
  wire  _T_2859 = _T_2839 ^ _T_2837; // @[AesSbox.scala 40:63]
  wire  _T_2861 = _T_2843 ^ _T_2853; // @[AesSbox.scala 40:63]
  wire  _T_2863 = _T_2855 ^ _T_2849; // @[AesSbox.scala 40:63]
  wire  _T_2865 = _T_2857 ^ _T_2853; // @[AesSbox.scala 40:63]
  wire  _T_2867 = _T_2859 ^ _T_2849; // @[AesSbox.scala 40:63]
  wire  _T_2869 = _T_2861 ^ _T_2823; // @[AesSbox.scala 40:63]
  wire  _T_2871 = _T_2867 ^ _T_2869; // @[AesSbox.scala 40:63]
  wire  _T_2873 = _T_2867 & _T_2863; // @[AesSbox.scala 41:63]
  wire  _T_2875 = _T_2865 ^ _T_2873; // @[AesSbox.scala 40:63]
  wire  _T_2877 = _T_2863 ^ _T_2865; // @[AesSbox.scala 40:63]
  wire  _T_2879 = _T_2869 ^ _T_2873; // @[AesSbox.scala 40:63]
  wire  _T_2881 = _T_2879 & _T_2877; // @[AesSbox.scala 41:63]
  wire  _T_2883 = _T_2875 & _T_2871; // @[AesSbox.scala 41:63]
  wire  _T_2885 = _T_2863 & _T_2869; // @[AesSbox.scala 41:63]
  wire  _T_2887 = _T_2877 & _T_2885; // @[AesSbox.scala 41:63]
  wire  _T_2889 = _T_2877 ^ _T_2873; // @[AesSbox.scala 40:63]
  wire  _T_2891 = _T_2865 & _T_2867; // @[AesSbox.scala 41:63]
  wire  _T_2893 = _T_2871 & _T_2891; // @[AesSbox.scala 41:63]
  wire  _T_2895 = _T_2871 ^ _T_2873; // @[AesSbox.scala 40:63]
  wire  _T_2897 = _T_2865 ^ _T_2881; // @[AesSbox.scala 40:63]
  wire  _T_2899 = _T_2887 ^ _T_2889; // @[AesSbox.scala 40:63]
  wire  _T_2901 = _T_2869 ^ _T_2883; // @[AesSbox.scala 40:63]
  wire  _T_2903 = _T_2893 ^ _T_2895; // @[AesSbox.scala 40:63]
  wire  _T_2905 = _T_2899 ^ _T_2903; // @[AesSbox.scala 40:63]
  wire  _T_2907 = _T_2897 ^ _T_2901; // @[AesSbox.scala 40:63]
  wire  _T_2909 = _T_2897 ^ _T_2899; // @[AesSbox.scala 40:63]
  wire  _T_2911 = _T_2901 ^ _T_2903; // @[AesSbox.scala 40:63]
  wire  _T_2913 = _T_2907 ^ _T_2905; // @[AesSbox.scala 40:63]
  wire  _T_2915 = _T_2911 & _T_2779; // @[AesSbox.scala 41:63]
  wire  _T_2917 = _T_2903 & _T_2791; // @[AesSbox.scala 41:63]
  wire  _T_2919 = _T_2901 & matrix_2_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_2921 = _T_2909 & _T_2811; // @[AesSbox.scala 41:63]
  wire  _T_2923 = _T_2899 & _T_2777; // @[AesSbox.scala 41:63]
  wire  _T_2925 = _T_2897 & _T_2803; // @[AesSbox.scala 41:63]
  wire  _T_2927 = _T_2907 & _T_2785; // @[AesSbox.scala 41:63]
  wire  _T_2929 = _T_2913 & _T_2815; // @[AesSbox.scala 41:63]
  wire  _T_2931 = _T_2905 & _T_2797; // @[AesSbox.scala 41:63]
  wire  _T_2933 = _T_2911 & _T_2807; // @[AesSbox.scala 41:63]
  wire  _T_2935 = _T_2903 & _T_2809; // @[AesSbox.scala 41:63]
  wire  _T_2937 = _T_2901 & _T_2789; // @[AesSbox.scala 41:63]
  wire  _T_2939 = _T_2909 & _T_2783; // @[AesSbox.scala 41:63]
  wire  _T_2941 = _T_2899 & _T_2787; // @[AesSbox.scala 41:63]
  wire  _T_2943 = _T_2897 & _T_2813; // @[AesSbox.scala 41:63]
  wire  _T_2945 = _T_2907 & _T_2773; // @[AesSbox.scala 41:63]
  wire  _T_2947 = _T_2913 & _T_2819; // @[AesSbox.scala 41:63]
  wire  _T_2949 = _T_2905 & _T_2801; // @[AesSbox.scala 41:63]
  wire  _T_2951 = _T_2945 ^ _T_2947; // @[AesSbox.scala 40:63]
  wire  _T_2953 = _T_2923 ^ _T_2935; // @[AesSbox.scala 40:63]
  wire  _T_2955 = _T_2929 ^ _T_2951; // @[AesSbox.scala 40:63]
  wire  _T_2957 = _T_2933 ^ _T_2953; // @[AesSbox.scala 40:63]
  wire  _T_2959 = _T_2919 ^ _T_2939; // @[AesSbox.scala 40:63]
  wire  _T_2961 = _T_2915 ^ _T_2921; // @[AesSbox.scala 40:63]
  wire  _T_2963 = _T_2951 ^ _T_2961; // @[AesSbox.scala 40:63]
  wire  _T_2965 = _T_2917 ^ _T_2957; // @[AesSbox.scala 40:63]
  wire  _T_2967 = _T_2915 ^ _T_2927; // @[AesSbox.scala 40:63]
  wire  _T_2969 = _T_2925 ^ _T_2941; // @[AesSbox.scala 40:63]
  wire  _T_2971 = _T_2931 ^ _T_2943; // @[AesSbox.scala 40:63]
  wire  _T_2973 = _T_2919 ^ _T_2965; // @[AesSbox.scala 40:63]
  wire  _T_2975 = _T_2959 ^ _T_2971; // @[AesSbox.scala 40:63]
  wire  _T_2977 = _T_2937 ^ _T_2953; // @[AesSbox.scala 40:63]
  wire  _T_2979 = _T_2921 ^ _T_2927; // @[AesSbox.scala 40:63]
  wire  _T_2981 = _T_2957 ^ _T_2979; // @[AesSbox.scala 40:63]
  wire  _T_2983 = _T_2949 ^ _T_2975; // @[AesSbox.scala 40:63]
  wire  _T_2985 = _T_2945 ^ _T_2967; // @[AesSbox.scala 40:63]
  wire  _T_2987 = _T_2959 ^ _T_2969; // @[AesSbox.scala 40:63]
  wire  _T_2988 = _T_2955 ^ _T_2981; // @[AesSbox.scala 40:63]
  wire  _T_2989 = _T_2983 ^ _T_2985; // @[AesSbox.scala 42:65]
  wire  _T_2990 = ~_T_2989; // @[AesSbox.scala 42:51]
  wire  _T_2992 = _T_2925 ^ _T_2951; // @[AesSbox.scala 40:63]
  wire  _T_2993 = _T_2963 ^ _T_2965; // @[AesSbox.scala 40:63]
  wire  _T_2994 = _T_2973 ^ _T_2992; // @[AesSbox.scala 40:63]
  wire  _T_2996 = _T_2923 ^ _T_2939; // @[AesSbox.scala 40:63]
  wire  _T_2998 = _T_2961 ^ _T_2977; // @[AesSbox.scala 40:63]
  wire  _T_2999 = _T_2963 ^ _T_2987; // @[AesSbox.scala 42:65]
  wire  _T_3000 = ~_T_2999; // @[AesSbox.scala 42:51]
  wire  _T_3002 = _T_2931 ^ _T_2969; // @[AesSbox.scala 40:63]
  wire  _T_3004 = _T_2996 ^ _T_3002; // @[AesSbox.scala 40:63]
  wire  _T_3006 = _T_2923 ^ _T_2967; // @[AesSbox.scala 40:63]
  wire  _T_3007 = _T_2955 ^ _T_3004; // @[AesSbox.scala 42:65]
  wire  _T_3008 = ~_T_3007; // @[AesSbox.scala 42:51]
  wire  _T_3010 = _T_2975 ^ _T_2998; // @[AesSbox.scala 40:63]
  wire  _T_3011 = _T_2955 ^ _T_3010; // @[AesSbox.scala 40:63]
  wire  _T_3013 = _T_2965 ^ _T_3006; // @[AesSbox.scala 40:63]
  wire  _T_3014 = _T_2955 ^ _T_3013; // @[AesSbox.scala 42:65]
  wire  _T_3015 = ~_T_3014; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_0_2 = {_T_2988,_T_3015,_T_2990,_T_2993,_T_2994,_T_3011,_T_3008,_T_3000}; // @[Cat.scala 29:58]
  wire  _T_3040 = matrix_2_3[1] ^ matrix_2_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_3042 = matrix_2_3[4] ^ matrix_2_3[7]; // @[AesSbox.scala 40:63]
  wire  _T_3044 = matrix_2_3[6] ^ matrix_2_3[5]; // @[AesSbox.scala 40:63]
  wire  _T_3046 = matrix_2_3[0] ^ _T_3044; // @[AesSbox.scala 40:63]
  wire  _T_3048 = _T_3040 ^ _T_3042; // @[AesSbox.scala 40:63]
  wire  _T_3050 = matrix_2_3[6] ^ matrix_2_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_3052 = matrix_2_3[7] ^ matrix_2_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_3054 = _T_3040 ^ _T_3050; // @[AesSbox.scala 40:63]
  wire  _T_3056 = matrix_2_3[1] ^ _T_3046; // @[AesSbox.scala 40:63]
  wire  _T_3058 = matrix_2_3[4] ^ _T_3046; // @[AesSbox.scala 40:63]
  wire  _T_3060 = matrix_2_3[0] ^ _T_3048; // @[AesSbox.scala 40:63]
  wire  _T_3062 = _T_3048 ^ _T_3050; // @[AesSbox.scala 40:63]
  wire  _T_3064 = matrix_2_3[5] ^ matrix_2_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_3066 = _T_3044 ^ _T_3048; // @[AesSbox.scala 40:63]
  wire  _T_3068 = matrix_2_3[2] ^ _T_3052; // @[AesSbox.scala 40:63]
  wire  _T_3070 = matrix_2_3[7] ^ matrix_2_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_3072 = matrix_2_3[0] ^ _T_3054; // @[AesSbox.scala 40:63]
  wire  _T_3074 = matrix_2_3[1] ^ matrix_2_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_3076 = _T_3042 ^ _T_3074; // @[AesSbox.scala 40:63]
  wire  _T_3078 = _T_3046 ^ _T_3068; // @[AesSbox.scala 40:63]
  wire  _T_3080 = _T_3040 ^ _T_3064; // @[AesSbox.scala 40:63]
  wire  _T_3082 = matrix_2_3[7] ^ _T_3046; // @[AesSbox.scala 40:63]
  wire  _T_3084 = _T_3080 ^ _T_3048; // @[AesSbox.scala 40:63]
  wire  _T_3086 = _T_3080 ^ _T_3052; // @[AesSbox.scala 40:63]
  wire  _T_3088 = _T_3052 ^ _T_3076; // @[AesSbox.scala 40:63]
  wire  _T_3090 = _T_3070 ^ _T_3066; // @[AesSbox.scala 40:63]
  wire  _T_3092 = _T_3082 ^ _T_3072; // @[AesSbox.scala 40:63]
  wire  _T_3094 = _T_3076 & _T_3048; // @[AesSbox.scala 41:63]
  wire  _T_3096 = _T_3078 & _T_3060; // @[AesSbox.scala 41:63]
  wire  _T_3098 = _T_3062 ^ _T_3094; // @[AesSbox.scala 40:63]
  wire  _T_3100 = _T_3058 & matrix_2_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_3102 = _T_3100 ^ _T_3094; // @[AesSbox.scala 40:63]
  wire  _T_3104 = _T_3052 & _T_3080; // @[AesSbox.scala 41:63]
  wire  _T_3106 = _T_3056 & _T_3046; // @[AesSbox.scala 41:63]
  wire  _T_3108 = _T_3086 ^ _T_3104; // @[AesSbox.scala 40:63]
  wire  _T_3110 = _T_3082 & _T_3072; // @[AesSbox.scala 41:63]
  wire  _T_3112 = _T_3110 ^ _T_3104; // @[AesSbox.scala 40:63]
  wire  _T_3114 = _T_3042 & _T_3054; // @[AesSbox.scala 41:63]
  wire  _T_3116 = _T_3088 & _T_3084; // @[AesSbox.scala 41:63]
  wire  _T_3118 = _T_3116 ^ _T_3114; // @[AesSbox.scala 40:63]
  wire  _T_3120 = _T_3070 & _T_3066; // @[AesSbox.scala 41:63]
  wire  _T_3122 = _T_3120 ^ _T_3114; // @[AesSbox.scala 40:63]
  wire  _T_3124 = _T_3098 ^ _T_3096; // @[AesSbox.scala 40:63]
  wire  _T_3126 = _T_3102 ^ _T_3090; // @[AesSbox.scala 40:63]
  wire  _T_3128 = _T_3108 ^ _T_3106; // @[AesSbox.scala 40:63]
  wire  _T_3130 = _T_3112 ^ _T_3122; // @[AesSbox.scala 40:63]
  wire  _T_3132 = _T_3124 ^ _T_3118; // @[AesSbox.scala 40:63]
  wire  _T_3134 = _T_3126 ^ _T_3122; // @[AesSbox.scala 40:63]
  wire  _T_3136 = _T_3128 ^ _T_3118; // @[AesSbox.scala 40:63]
  wire  _T_3138 = _T_3130 ^ _T_3092; // @[AesSbox.scala 40:63]
  wire  _T_3140 = _T_3136 ^ _T_3138; // @[AesSbox.scala 40:63]
  wire  _T_3142 = _T_3136 & _T_3132; // @[AesSbox.scala 41:63]
  wire  _T_3144 = _T_3134 ^ _T_3142; // @[AesSbox.scala 40:63]
  wire  _T_3146 = _T_3132 ^ _T_3134; // @[AesSbox.scala 40:63]
  wire  _T_3148 = _T_3138 ^ _T_3142; // @[AesSbox.scala 40:63]
  wire  _T_3150 = _T_3148 & _T_3146; // @[AesSbox.scala 41:63]
  wire  _T_3152 = _T_3144 & _T_3140; // @[AesSbox.scala 41:63]
  wire  _T_3154 = _T_3132 & _T_3138; // @[AesSbox.scala 41:63]
  wire  _T_3156 = _T_3146 & _T_3154; // @[AesSbox.scala 41:63]
  wire  _T_3158 = _T_3146 ^ _T_3142; // @[AesSbox.scala 40:63]
  wire  _T_3160 = _T_3134 & _T_3136; // @[AesSbox.scala 41:63]
  wire  _T_3162 = _T_3140 & _T_3160; // @[AesSbox.scala 41:63]
  wire  _T_3164 = _T_3140 ^ _T_3142; // @[AesSbox.scala 40:63]
  wire  _T_3166 = _T_3134 ^ _T_3150; // @[AesSbox.scala 40:63]
  wire  _T_3168 = _T_3156 ^ _T_3158; // @[AesSbox.scala 40:63]
  wire  _T_3170 = _T_3138 ^ _T_3152; // @[AesSbox.scala 40:63]
  wire  _T_3172 = _T_3162 ^ _T_3164; // @[AesSbox.scala 40:63]
  wire  _T_3174 = _T_3168 ^ _T_3172; // @[AesSbox.scala 40:63]
  wire  _T_3176 = _T_3166 ^ _T_3170; // @[AesSbox.scala 40:63]
  wire  _T_3178 = _T_3166 ^ _T_3168; // @[AesSbox.scala 40:63]
  wire  _T_3180 = _T_3170 ^ _T_3172; // @[AesSbox.scala 40:63]
  wire  _T_3182 = _T_3176 ^ _T_3174; // @[AesSbox.scala 40:63]
  wire  _T_3184 = _T_3180 & _T_3048; // @[AesSbox.scala 41:63]
  wire  _T_3186 = _T_3172 & _T_3060; // @[AesSbox.scala 41:63]
  wire  _T_3188 = _T_3170 & matrix_2_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_3190 = _T_3178 & _T_3080; // @[AesSbox.scala 41:63]
  wire  _T_3192 = _T_3168 & _T_3046; // @[AesSbox.scala 41:63]
  wire  _T_3194 = _T_3166 & _T_3072; // @[AesSbox.scala 41:63]
  wire  _T_3196 = _T_3176 & _T_3054; // @[AesSbox.scala 41:63]
  wire  _T_3198 = _T_3182 & _T_3084; // @[AesSbox.scala 41:63]
  wire  _T_3200 = _T_3174 & _T_3066; // @[AesSbox.scala 41:63]
  wire  _T_3202 = _T_3180 & _T_3076; // @[AesSbox.scala 41:63]
  wire  _T_3204 = _T_3172 & _T_3078; // @[AesSbox.scala 41:63]
  wire  _T_3206 = _T_3170 & _T_3058; // @[AesSbox.scala 41:63]
  wire  _T_3208 = _T_3178 & _T_3052; // @[AesSbox.scala 41:63]
  wire  _T_3210 = _T_3168 & _T_3056; // @[AesSbox.scala 41:63]
  wire  _T_3212 = _T_3166 & _T_3082; // @[AesSbox.scala 41:63]
  wire  _T_3214 = _T_3176 & _T_3042; // @[AesSbox.scala 41:63]
  wire  _T_3216 = _T_3182 & _T_3088; // @[AesSbox.scala 41:63]
  wire  _T_3218 = _T_3174 & _T_3070; // @[AesSbox.scala 41:63]
  wire  _T_3220 = _T_3214 ^ _T_3216; // @[AesSbox.scala 40:63]
  wire  _T_3222 = _T_3192 ^ _T_3204; // @[AesSbox.scala 40:63]
  wire  _T_3224 = _T_3198 ^ _T_3220; // @[AesSbox.scala 40:63]
  wire  _T_3226 = _T_3202 ^ _T_3222; // @[AesSbox.scala 40:63]
  wire  _T_3228 = _T_3188 ^ _T_3208; // @[AesSbox.scala 40:63]
  wire  _T_3230 = _T_3184 ^ _T_3190; // @[AesSbox.scala 40:63]
  wire  _T_3232 = _T_3220 ^ _T_3230; // @[AesSbox.scala 40:63]
  wire  _T_3234 = _T_3186 ^ _T_3226; // @[AesSbox.scala 40:63]
  wire  _T_3236 = _T_3184 ^ _T_3196; // @[AesSbox.scala 40:63]
  wire  _T_3238 = _T_3194 ^ _T_3210; // @[AesSbox.scala 40:63]
  wire  _T_3240 = _T_3200 ^ _T_3212; // @[AesSbox.scala 40:63]
  wire  _T_3242 = _T_3188 ^ _T_3234; // @[AesSbox.scala 40:63]
  wire  _T_3244 = _T_3228 ^ _T_3240; // @[AesSbox.scala 40:63]
  wire  _T_3246 = _T_3206 ^ _T_3222; // @[AesSbox.scala 40:63]
  wire  _T_3248 = _T_3190 ^ _T_3196; // @[AesSbox.scala 40:63]
  wire  _T_3250 = _T_3226 ^ _T_3248; // @[AesSbox.scala 40:63]
  wire  _T_3252 = _T_3218 ^ _T_3244; // @[AesSbox.scala 40:63]
  wire  _T_3254 = _T_3214 ^ _T_3236; // @[AesSbox.scala 40:63]
  wire  _T_3256 = _T_3228 ^ _T_3238; // @[AesSbox.scala 40:63]
  wire  _T_3257 = _T_3224 ^ _T_3250; // @[AesSbox.scala 40:63]
  wire  _T_3258 = _T_3252 ^ _T_3254; // @[AesSbox.scala 42:65]
  wire  _T_3259 = ~_T_3258; // @[AesSbox.scala 42:51]
  wire  _T_3261 = _T_3194 ^ _T_3220; // @[AesSbox.scala 40:63]
  wire  _T_3262 = _T_3232 ^ _T_3234; // @[AesSbox.scala 40:63]
  wire  _T_3263 = _T_3242 ^ _T_3261; // @[AesSbox.scala 40:63]
  wire  _T_3265 = _T_3192 ^ _T_3208; // @[AesSbox.scala 40:63]
  wire  _T_3267 = _T_3230 ^ _T_3246; // @[AesSbox.scala 40:63]
  wire  _T_3268 = _T_3232 ^ _T_3256; // @[AesSbox.scala 42:65]
  wire  _T_3269 = ~_T_3268; // @[AesSbox.scala 42:51]
  wire  _T_3271 = _T_3200 ^ _T_3238; // @[AesSbox.scala 40:63]
  wire  _T_3273 = _T_3265 ^ _T_3271; // @[AesSbox.scala 40:63]
  wire  _T_3275 = _T_3192 ^ _T_3236; // @[AesSbox.scala 40:63]
  wire  _T_3276 = _T_3224 ^ _T_3273; // @[AesSbox.scala 42:65]
  wire  _T_3277 = ~_T_3276; // @[AesSbox.scala 42:51]
  wire  _T_3279 = _T_3244 ^ _T_3267; // @[AesSbox.scala 40:63]
  wire  _T_3280 = _T_3224 ^ _T_3279; // @[AesSbox.scala 40:63]
  wire  _T_3282 = _T_3234 ^ _T_3275; // @[AesSbox.scala 40:63]
  wire  _T_3283 = _T_3224 ^ _T_3282; // @[AesSbox.scala 42:65]
  wire  _T_3284 = ~_T_3283; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_3_3 = {_T_3257,_T_3284,_T_3259,_T_3262,_T_3263,_T_3280,_T_3277,_T_3269}; // @[Cat.scala 29:58]
  wire  _T_3310 = matrix_3_0[1] ^ matrix_3_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_3312 = matrix_3_0[4] ^ matrix_3_0[7]; // @[AesSbox.scala 40:63]
  wire  _T_3314 = matrix_3_0[6] ^ matrix_3_0[5]; // @[AesSbox.scala 40:63]
  wire  _T_3316 = matrix_3_0[0] ^ _T_3314; // @[AesSbox.scala 40:63]
  wire  _T_3318 = _T_3310 ^ _T_3312; // @[AesSbox.scala 40:63]
  wire  _T_3320 = matrix_3_0[6] ^ matrix_3_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_3322 = matrix_3_0[7] ^ matrix_3_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_3324 = _T_3310 ^ _T_3320; // @[AesSbox.scala 40:63]
  wire  _T_3326 = matrix_3_0[1] ^ _T_3316; // @[AesSbox.scala 40:63]
  wire  _T_3328 = matrix_3_0[4] ^ _T_3316; // @[AesSbox.scala 40:63]
  wire  _T_3330 = matrix_3_0[0] ^ _T_3318; // @[AesSbox.scala 40:63]
  wire  _T_3332 = _T_3318 ^ _T_3320; // @[AesSbox.scala 40:63]
  wire  _T_3334 = matrix_3_0[5] ^ matrix_3_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_3336 = _T_3314 ^ _T_3318; // @[AesSbox.scala 40:63]
  wire  _T_3338 = matrix_3_0[2] ^ _T_3322; // @[AesSbox.scala 40:63]
  wire  _T_3340 = matrix_3_0[7] ^ matrix_3_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_3342 = matrix_3_0[0] ^ _T_3324; // @[AesSbox.scala 40:63]
  wire  _T_3344 = matrix_3_0[1] ^ matrix_3_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_3346 = _T_3312 ^ _T_3344; // @[AesSbox.scala 40:63]
  wire  _T_3348 = _T_3316 ^ _T_3338; // @[AesSbox.scala 40:63]
  wire  _T_3350 = _T_3310 ^ _T_3334; // @[AesSbox.scala 40:63]
  wire  _T_3352 = matrix_3_0[7] ^ _T_3316; // @[AesSbox.scala 40:63]
  wire  _T_3354 = _T_3350 ^ _T_3318; // @[AesSbox.scala 40:63]
  wire  _T_3356 = _T_3350 ^ _T_3322; // @[AesSbox.scala 40:63]
  wire  _T_3358 = _T_3322 ^ _T_3346; // @[AesSbox.scala 40:63]
  wire  _T_3360 = _T_3340 ^ _T_3336; // @[AesSbox.scala 40:63]
  wire  _T_3362 = _T_3352 ^ _T_3342; // @[AesSbox.scala 40:63]
  wire  _T_3364 = _T_3346 & _T_3318; // @[AesSbox.scala 41:63]
  wire  _T_3366 = _T_3348 & _T_3330; // @[AesSbox.scala 41:63]
  wire  _T_3368 = _T_3332 ^ _T_3364; // @[AesSbox.scala 40:63]
  wire  _T_3370 = _T_3328 & matrix_3_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_3372 = _T_3370 ^ _T_3364; // @[AesSbox.scala 40:63]
  wire  _T_3374 = _T_3322 & _T_3350; // @[AesSbox.scala 41:63]
  wire  _T_3376 = _T_3326 & _T_3316; // @[AesSbox.scala 41:63]
  wire  _T_3378 = _T_3356 ^ _T_3374; // @[AesSbox.scala 40:63]
  wire  _T_3380 = _T_3352 & _T_3342; // @[AesSbox.scala 41:63]
  wire  _T_3382 = _T_3380 ^ _T_3374; // @[AesSbox.scala 40:63]
  wire  _T_3384 = _T_3312 & _T_3324; // @[AesSbox.scala 41:63]
  wire  _T_3386 = _T_3358 & _T_3354; // @[AesSbox.scala 41:63]
  wire  _T_3388 = _T_3386 ^ _T_3384; // @[AesSbox.scala 40:63]
  wire  _T_3390 = _T_3340 & _T_3336; // @[AesSbox.scala 41:63]
  wire  _T_3392 = _T_3390 ^ _T_3384; // @[AesSbox.scala 40:63]
  wire  _T_3394 = _T_3368 ^ _T_3366; // @[AesSbox.scala 40:63]
  wire  _T_3396 = _T_3372 ^ _T_3360; // @[AesSbox.scala 40:63]
  wire  _T_3398 = _T_3378 ^ _T_3376; // @[AesSbox.scala 40:63]
  wire  _T_3400 = _T_3382 ^ _T_3392; // @[AesSbox.scala 40:63]
  wire  _T_3402 = _T_3394 ^ _T_3388; // @[AesSbox.scala 40:63]
  wire  _T_3404 = _T_3396 ^ _T_3392; // @[AesSbox.scala 40:63]
  wire  _T_3406 = _T_3398 ^ _T_3388; // @[AesSbox.scala 40:63]
  wire  _T_3408 = _T_3400 ^ _T_3362; // @[AesSbox.scala 40:63]
  wire  _T_3410 = _T_3406 ^ _T_3408; // @[AesSbox.scala 40:63]
  wire  _T_3412 = _T_3406 & _T_3402; // @[AesSbox.scala 41:63]
  wire  _T_3414 = _T_3404 ^ _T_3412; // @[AesSbox.scala 40:63]
  wire  _T_3416 = _T_3402 ^ _T_3404; // @[AesSbox.scala 40:63]
  wire  _T_3418 = _T_3408 ^ _T_3412; // @[AesSbox.scala 40:63]
  wire  _T_3420 = _T_3418 & _T_3416; // @[AesSbox.scala 41:63]
  wire  _T_3422 = _T_3414 & _T_3410; // @[AesSbox.scala 41:63]
  wire  _T_3424 = _T_3402 & _T_3408; // @[AesSbox.scala 41:63]
  wire  _T_3426 = _T_3416 & _T_3424; // @[AesSbox.scala 41:63]
  wire  _T_3428 = _T_3416 ^ _T_3412; // @[AesSbox.scala 40:63]
  wire  _T_3430 = _T_3404 & _T_3406; // @[AesSbox.scala 41:63]
  wire  _T_3432 = _T_3410 & _T_3430; // @[AesSbox.scala 41:63]
  wire  _T_3434 = _T_3410 ^ _T_3412; // @[AesSbox.scala 40:63]
  wire  _T_3436 = _T_3404 ^ _T_3420; // @[AesSbox.scala 40:63]
  wire  _T_3438 = _T_3426 ^ _T_3428; // @[AesSbox.scala 40:63]
  wire  _T_3440 = _T_3408 ^ _T_3422; // @[AesSbox.scala 40:63]
  wire  _T_3442 = _T_3432 ^ _T_3434; // @[AesSbox.scala 40:63]
  wire  _T_3444 = _T_3438 ^ _T_3442; // @[AesSbox.scala 40:63]
  wire  _T_3446 = _T_3436 ^ _T_3440; // @[AesSbox.scala 40:63]
  wire  _T_3448 = _T_3436 ^ _T_3438; // @[AesSbox.scala 40:63]
  wire  _T_3450 = _T_3440 ^ _T_3442; // @[AesSbox.scala 40:63]
  wire  _T_3452 = _T_3446 ^ _T_3444; // @[AesSbox.scala 40:63]
  wire  _T_3454 = _T_3450 & _T_3318; // @[AesSbox.scala 41:63]
  wire  _T_3456 = _T_3442 & _T_3330; // @[AesSbox.scala 41:63]
  wire  _T_3458 = _T_3440 & matrix_3_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_3460 = _T_3448 & _T_3350; // @[AesSbox.scala 41:63]
  wire  _T_3462 = _T_3438 & _T_3316; // @[AesSbox.scala 41:63]
  wire  _T_3464 = _T_3436 & _T_3342; // @[AesSbox.scala 41:63]
  wire  _T_3466 = _T_3446 & _T_3324; // @[AesSbox.scala 41:63]
  wire  _T_3468 = _T_3452 & _T_3354; // @[AesSbox.scala 41:63]
  wire  _T_3470 = _T_3444 & _T_3336; // @[AesSbox.scala 41:63]
  wire  _T_3472 = _T_3450 & _T_3346; // @[AesSbox.scala 41:63]
  wire  _T_3474 = _T_3442 & _T_3348; // @[AesSbox.scala 41:63]
  wire  _T_3476 = _T_3440 & _T_3328; // @[AesSbox.scala 41:63]
  wire  _T_3478 = _T_3448 & _T_3322; // @[AesSbox.scala 41:63]
  wire  _T_3480 = _T_3438 & _T_3326; // @[AesSbox.scala 41:63]
  wire  _T_3482 = _T_3436 & _T_3352; // @[AesSbox.scala 41:63]
  wire  _T_3484 = _T_3446 & _T_3312; // @[AesSbox.scala 41:63]
  wire  _T_3486 = _T_3452 & _T_3358; // @[AesSbox.scala 41:63]
  wire  _T_3488 = _T_3444 & _T_3340; // @[AesSbox.scala 41:63]
  wire  _T_3490 = _T_3484 ^ _T_3486; // @[AesSbox.scala 40:63]
  wire  _T_3492 = _T_3462 ^ _T_3474; // @[AesSbox.scala 40:63]
  wire  _T_3494 = _T_3468 ^ _T_3490; // @[AesSbox.scala 40:63]
  wire  _T_3496 = _T_3472 ^ _T_3492; // @[AesSbox.scala 40:63]
  wire  _T_3498 = _T_3458 ^ _T_3478; // @[AesSbox.scala 40:63]
  wire  _T_3500 = _T_3454 ^ _T_3460; // @[AesSbox.scala 40:63]
  wire  _T_3502 = _T_3490 ^ _T_3500; // @[AesSbox.scala 40:63]
  wire  _T_3504 = _T_3456 ^ _T_3496; // @[AesSbox.scala 40:63]
  wire  _T_3506 = _T_3454 ^ _T_3466; // @[AesSbox.scala 40:63]
  wire  _T_3508 = _T_3464 ^ _T_3480; // @[AesSbox.scala 40:63]
  wire  _T_3510 = _T_3470 ^ _T_3482; // @[AesSbox.scala 40:63]
  wire  _T_3512 = _T_3458 ^ _T_3504; // @[AesSbox.scala 40:63]
  wire  _T_3514 = _T_3498 ^ _T_3510; // @[AesSbox.scala 40:63]
  wire  _T_3516 = _T_3476 ^ _T_3492; // @[AesSbox.scala 40:63]
  wire  _T_3518 = _T_3460 ^ _T_3466; // @[AesSbox.scala 40:63]
  wire  _T_3520 = _T_3496 ^ _T_3518; // @[AesSbox.scala 40:63]
  wire  _T_3522 = _T_3488 ^ _T_3514; // @[AesSbox.scala 40:63]
  wire  _T_3524 = _T_3484 ^ _T_3506; // @[AesSbox.scala 40:63]
  wire  _T_3526 = _T_3498 ^ _T_3508; // @[AesSbox.scala 40:63]
  wire  _T_3527 = _T_3494 ^ _T_3520; // @[AesSbox.scala 40:63]
  wire  _T_3528 = _T_3522 ^ _T_3524; // @[AesSbox.scala 42:65]
  wire  _T_3529 = ~_T_3528; // @[AesSbox.scala 42:51]
  wire  _T_3531 = _T_3464 ^ _T_3490; // @[AesSbox.scala 40:63]
  wire  _T_3532 = _T_3502 ^ _T_3504; // @[AesSbox.scala 40:63]
  wire  _T_3533 = _T_3512 ^ _T_3531; // @[AesSbox.scala 40:63]
  wire  _T_3535 = _T_3462 ^ _T_3478; // @[AesSbox.scala 40:63]
  wire  _T_3537 = _T_3500 ^ _T_3516; // @[AesSbox.scala 40:63]
  wire  _T_3538 = _T_3502 ^ _T_3526; // @[AesSbox.scala 42:65]
  wire  _T_3539 = ~_T_3538; // @[AesSbox.scala 42:51]
  wire  _T_3541 = _T_3470 ^ _T_3508; // @[AesSbox.scala 40:63]
  wire  _T_3543 = _T_3535 ^ _T_3541; // @[AesSbox.scala 40:63]
  wire  _T_3545 = _T_3462 ^ _T_3506; // @[AesSbox.scala 40:63]
  wire  _T_3546 = _T_3494 ^ _T_3543; // @[AesSbox.scala 42:65]
  wire  _T_3547 = ~_T_3546; // @[AesSbox.scala 42:51]
  wire  _T_3549 = _T_3514 ^ _T_3537; // @[AesSbox.scala 40:63]
  wire  _T_3550 = _T_3494 ^ _T_3549; // @[AesSbox.scala 40:63]
  wire  _T_3552 = _T_3504 ^ _T_3545; // @[AesSbox.scala 40:63]
  wire  _T_3553 = _T_3494 ^ _T_3552; // @[AesSbox.scala 42:65]
  wire  _T_3554 = ~_T_3553; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_3_0 = {_T_3527,_T_3554,_T_3529,_T_3532,_T_3533,_T_3550,_T_3547,_T_3539}; // @[Cat.scala 29:58]
  wire  _T_3579 = matrix_3_1[1] ^ matrix_3_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_3581 = matrix_3_1[4] ^ matrix_3_1[7]; // @[AesSbox.scala 40:63]
  wire  _T_3583 = matrix_3_1[6] ^ matrix_3_1[5]; // @[AesSbox.scala 40:63]
  wire  _T_3585 = matrix_3_1[0] ^ _T_3583; // @[AesSbox.scala 40:63]
  wire  _T_3587 = _T_3579 ^ _T_3581; // @[AesSbox.scala 40:63]
  wire  _T_3589 = matrix_3_1[6] ^ matrix_3_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_3591 = matrix_3_1[7] ^ matrix_3_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_3593 = _T_3579 ^ _T_3589; // @[AesSbox.scala 40:63]
  wire  _T_3595 = matrix_3_1[1] ^ _T_3585; // @[AesSbox.scala 40:63]
  wire  _T_3597 = matrix_3_1[4] ^ _T_3585; // @[AesSbox.scala 40:63]
  wire  _T_3599 = matrix_3_1[0] ^ _T_3587; // @[AesSbox.scala 40:63]
  wire  _T_3601 = _T_3587 ^ _T_3589; // @[AesSbox.scala 40:63]
  wire  _T_3603 = matrix_3_1[5] ^ matrix_3_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_3605 = _T_3583 ^ _T_3587; // @[AesSbox.scala 40:63]
  wire  _T_3607 = matrix_3_1[2] ^ _T_3591; // @[AesSbox.scala 40:63]
  wire  _T_3609 = matrix_3_1[7] ^ matrix_3_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_3611 = matrix_3_1[0] ^ _T_3593; // @[AesSbox.scala 40:63]
  wire  _T_3613 = matrix_3_1[1] ^ matrix_3_1[2]; // @[AesSbox.scala 40:63]
  wire  _T_3615 = _T_3581 ^ _T_3613; // @[AesSbox.scala 40:63]
  wire  _T_3617 = _T_3585 ^ _T_3607; // @[AesSbox.scala 40:63]
  wire  _T_3619 = _T_3579 ^ _T_3603; // @[AesSbox.scala 40:63]
  wire  _T_3621 = matrix_3_1[7] ^ _T_3585; // @[AesSbox.scala 40:63]
  wire  _T_3623 = _T_3619 ^ _T_3587; // @[AesSbox.scala 40:63]
  wire  _T_3625 = _T_3619 ^ _T_3591; // @[AesSbox.scala 40:63]
  wire  _T_3627 = _T_3591 ^ _T_3615; // @[AesSbox.scala 40:63]
  wire  _T_3629 = _T_3609 ^ _T_3605; // @[AesSbox.scala 40:63]
  wire  _T_3631 = _T_3621 ^ _T_3611; // @[AesSbox.scala 40:63]
  wire  _T_3633 = _T_3615 & _T_3587; // @[AesSbox.scala 41:63]
  wire  _T_3635 = _T_3617 & _T_3599; // @[AesSbox.scala 41:63]
  wire  _T_3637 = _T_3601 ^ _T_3633; // @[AesSbox.scala 40:63]
  wire  _T_3639 = _T_3597 & matrix_3_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_3641 = _T_3639 ^ _T_3633; // @[AesSbox.scala 40:63]
  wire  _T_3643 = _T_3591 & _T_3619; // @[AesSbox.scala 41:63]
  wire  _T_3645 = _T_3595 & _T_3585; // @[AesSbox.scala 41:63]
  wire  _T_3647 = _T_3625 ^ _T_3643; // @[AesSbox.scala 40:63]
  wire  _T_3649 = _T_3621 & _T_3611; // @[AesSbox.scala 41:63]
  wire  _T_3651 = _T_3649 ^ _T_3643; // @[AesSbox.scala 40:63]
  wire  _T_3653 = _T_3581 & _T_3593; // @[AesSbox.scala 41:63]
  wire  _T_3655 = _T_3627 & _T_3623; // @[AesSbox.scala 41:63]
  wire  _T_3657 = _T_3655 ^ _T_3653; // @[AesSbox.scala 40:63]
  wire  _T_3659 = _T_3609 & _T_3605; // @[AesSbox.scala 41:63]
  wire  _T_3661 = _T_3659 ^ _T_3653; // @[AesSbox.scala 40:63]
  wire  _T_3663 = _T_3637 ^ _T_3635; // @[AesSbox.scala 40:63]
  wire  _T_3665 = _T_3641 ^ _T_3629; // @[AesSbox.scala 40:63]
  wire  _T_3667 = _T_3647 ^ _T_3645; // @[AesSbox.scala 40:63]
  wire  _T_3669 = _T_3651 ^ _T_3661; // @[AesSbox.scala 40:63]
  wire  _T_3671 = _T_3663 ^ _T_3657; // @[AesSbox.scala 40:63]
  wire  _T_3673 = _T_3665 ^ _T_3661; // @[AesSbox.scala 40:63]
  wire  _T_3675 = _T_3667 ^ _T_3657; // @[AesSbox.scala 40:63]
  wire  _T_3677 = _T_3669 ^ _T_3631; // @[AesSbox.scala 40:63]
  wire  _T_3679 = _T_3675 ^ _T_3677; // @[AesSbox.scala 40:63]
  wire  _T_3681 = _T_3675 & _T_3671; // @[AesSbox.scala 41:63]
  wire  _T_3683 = _T_3673 ^ _T_3681; // @[AesSbox.scala 40:63]
  wire  _T_3685 = _T_3671 ^ _T_3673; // @[AesSbox.scala 40:63]
  wire  _T_3687 = _T_3677 ^ _T_3681; // @[AesSbox.scala 40:63]
  wire  _T_3689 = _T_3687 & _T_3685; // @[AesSbox.scala 41:63]
  wire  _T_3691 = _T_3683 & _T_3679; // @[AesSbox.scala 41:63]
  wire  _T_3693 = _T_3671 & _T_3677; // @[AesSbox.scala 41:63]
  wire  _T_3695 = _T_3685 & _T_3693; // @[AesSbox.scala 41:63]
  wire  _T_3697 = _T_3685 ^ _T_3681; // @[AesSbox.scala 40:63]
  wire  _T_3699 = _T_3673 & _T_3675; // @[AesSbox.scala 41:63]
  wire  _T_3701 = _T_3679 & _T_3699; // @[AesSbox.scala 41:63]
  wire  _T_3703 = _T_3679 ^ _T_3681; // @[AesSbox.scala 40:63]
  wire  _T_3705 = _T_3673 ^ _T_3689; // @[AesSbox.scala 40:63]
  wire  _T_3707 = _T_3695 ^ _T_3697; // @[AesSbox.scala 40:63]
  wire  _T_3709 = _T_3677 ^ _T_3691; // @[AesSbox.scala 40:63]
  wire  _T_3711 = _T_3701 ^ _T_3703; // @[AesSbox.scala 40:63]
  wire  _T_3713 = _T_3707 ^ _T_3711; // @[AesSbox.scala 40:63]
  wire  _T_3715 = _T_3705 ^ _T_3709; // @[AesSbox.scala 40:63]
  wire  _T_3717 = _T_3705 ^ _T_3707; // @[AesSbox.scala 40:63]
  wire  _T_3719 = _T_3709 ^ _T_3711; // @[AesSbox.scala 40:63]
  wire  _T_3721 = _T_3715 ^ _T_3713; // @[AesSbox.scala 40:63]
  wire  _T_3723 = _T_3719 & _T_3587; // @[AesSbox.scala 41:63]
  wire  _T_3725 = _T_3711 & _T_3599; // @[AesSbox.scala 41:63]
  wire  _T_3727 = _T_3709 & matrix_3_1[0]; // @[AesSbox.scala 41:63]
  wire  _T_3729 = _T_3717 & _T_3619; // @[AesSbox.scala 41:63]
  wire  _T_3731 = _T_3707 & _T_3585; // @[AesSbox.scala 41:63]
  wire  _T_3733 = _T_3705 & _T_3611; // @[AesSbox.scala 41:63]
  wire  _T_3735 = _T_3715 & _T_3593; // @[AesSbox.scala 41:63]
  wire  _T_3737 = _T_3721 & _T_3623; // @[AesSbox.scala 41:63]
  wire  _T_3739 = _T_3713 & _T_3605; // @[AesSbox.scala 41:63]
  wire  _T_3741 = _T_3719 & _T_3615; // @[AesSbox.scala 41:63]
  wire  _T_3743 = _T_3711 & _T_3617; // @[AesSbox.scala 41:63]
  wire  _T_3745 = _T_3709 & _T_3597; // @[AesSbox.scala 41:63]
  wire  _T_3747 = _T_3717 & _T_3591; // @[AesSbox.scala 41:63]
  wire  _T_3749 = _T_3707 & _T_3595; // @[AesSbox.scala 41:63]
  wire  _T_3751 = _T_3705 & _T_3621; // @[AesSbox.scala 41:63]
  wire  _T_3753 = _T_3715 & _T_3581; // @[AesSbox.scala 41:63]
  wire  _T_3755 = _T_3721 & _T_3627; // @[AesSbox.scala 41:63]
  wire  _T_3757 = _T_3713 & _T_3609; // @[AesSbox.scala 41:63]
  wire  _T_3759 = _T_3753 ^ _T_3755; // @[AesSbox.scala 40:63]
  wire  _T_3761 = _T_3731 ^ _T_3743; // @[AesSbox.scala 40:63]
  wire  _T_3763 = _T_3737 ^ _T_3759; // @[AesSbox.scala 40:63]
  wire  _T_3765 = _T_3741 ^ _T_3761; // @[AesSbox.scala 40:63]
  wire  _T_3767 = _T_3727 ^ _T_3747; // @[AesSbox.scala 40:63]
  wire  _T_3769 = _T_3723 ^ _T_3729; // @[AesSbox.scala 40:63]
  wire  _T_3771 = _T_3759 ^ _T_3769; // @[AesSbox.scala 40:63]
  wire  _T_3773 = _T_3725 ^ _T_3765; // @[AesSbox.scala 40:63]
  wire  _T_3775 = _T_3723 ^ _T_3735; // @[AesSbox.scala 40:63]
  wire  _T_3777 = _T_3733 ^ _T_3749; // @[AesSbox.scala 40:63]
  wire  _T_3779 = _T_3739 ^ _T_3751; // @[AesSbox.scala 40:63]
  wire  _T_3781 = _T_3727 ^ _T_3773; // @[AesSbox.scala 40:63]
  wire  _T_3783 = _T_3767 ^ _T_3779; // @[AesSbox.scala 40:63]
  wire  _T_3785 = _T_3745 ^ _T_3761; // @[AesSbox.scala 40:63]
  wire  _T_3787 = _T_3729 ^ _T_3735; // @[AesSbox.scala 40:63]
  wire  _T_3789 = _T_3765 ^ _T_3787; // @[AesSbox.scala 40:63]
  wire  _T_3791 = _T_3757 ^ _T_3783; // @[AesSbox.scala 40:63]
  wire  _T_3793 = _T_3753 ^ _T_3775; // @[AesSbox.scala 40:63]
  wire  _T_3795 = _T_3767 ^ _T_3777; // @[AesSbox.scala 40:63]
  wire  _T_3796 = _T_3763 ^ _T_3789; // @[AesSbox.scala 40:63]
  wire  _T_3797 = _T_3791 ^ _T_3793; // @[AesSbox.scala 42:65]
  wire  _T_3798 = ~_T_3797; // @[AesSbox.scala 42:51]
  wire  _T_3800 = _T_3733 ^ _T_3759; // @[AesSbox.scala 40:63]
  wire  _T_3801 = _T_3771 ^ _T_3773; // @[AesSbox.scala 40:63]
  wire  _T_3802 = _T_3781 ^ _T_3800; // @[AesSbox.scala 40:63]
  wire  _T_3804 = _T_3731 ^ _T_3747; // @[AesSbox.scala 40:63]
  wire  _T_3806 = _T_3769 ^ _T_3785; // @[AesSbox.scala 40:63]
  wire  _T_3807 = _T_3771 ^ _T_3795; // @[AesSbox.scala 42:65]
  wire  _T_3808 = ~_T_3807; // @[AesSbox.scala 42:51]
  wire  _T_3810 = _T_3739 ^ _T_3777; // @[AesSbox.scala 40:63]
  wire  _T_3812 = _T_3804 ^ _T_3810; // @[AesSbox.scala 40:63]
  wire  _T_3814 = _T_3731 ^ _T_3775; // @[AesSbox.scala 40:63]
  wire  _T_3815 = _T_3763 ^ _T_3812; // @[AesSbox.scala 42:65]
  wire  _T_3816 = ~_T_3815; // @[AesSbox.scala 42:51]
  wire  _T_3818 = _T_3783 ^ _T_3806; // @[AesSbox.scala 40:63]
  wire  _T_3819 = _T_3763 ^ _T_3818; // @[AesSbox.scala 40:63]
  wire  _T_3821 = _T_3773 ^ _T_3814; // @[AesSbox.scala 40:63]
  wire  _T_3822 = _T_3763 ^ _T_3821; // @[AesSbox.scala 42:65]
  wire  _T_3823 = ~_T_3822; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_2_1 = {_T_3796,_T_3823,_T_3798,_T_3801,_T_3802,_T_3819,_T_3816,_T_3808}; // @[Cat.scala 29:58]
  wire  _T_3848 = matrix_3_2[1] ^ matrix_3_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_3850 = matrix_3_2[4] ^ matrix_3_2[7]; // @[AesSbox.scala 40:63]
  wire  _T_3852 = matrix_3_2[6] ^ matrix_3_2[5]; // @[AesSbox.scala 40:63]
  wire  _T_3854 = matrix_3_2[0] ^ _T_3852; // @[AesSbox.scala 40:63]
  wire  _T_3856 = _T_3848 ^ _T_3850; // @[AesSbox.scala 40:63]
  wire  _T_3858 = matrix_3_2[6] ^ matrix_3_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_3860 = matrix_3_2[7] ^ matrix_3_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_3862 = _T_3848 ^ _T_3858; // @[AesSbox.scala 40:63]
  wire  _T_3864 = matrix_3_2[1] ^ _T_3854; // @[AesSbox.scala 40:63]
  wire  _T_3866 = matrix_3_2[4] ^ _T_3854; // @[AesSbox.scala 40:63]
  wire  _T_3868 = matrix_3_2[0] ^ _T_3856; // @[AesSbox.scala 40:63]
  wire  _T_3870 = _T_3856 ^ _T_3858; // @[AesSbox.scala 40:63]
  wire  _T_3872 = matrix_3_2[5] ^ matrix_3_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_3874 = _T_3852 ^ _T_3856; // @[AesSbox.scala 40:63]
  wire  _T_3876 = matrix_3_2[2] ^ _T_3860; // @[AesSbox.scala 40:63]
  wire  _T_3878 = matrix_3_2[7] ^ matrix_3_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_3880 = matrix_3_2[0] ^ _T_3862; // @[AesSbox.scala 40:63]
  wire  _T_3882 = matrix_3_2[1] ^ matrix_3_2[2]; // @[AesSbox.scala 40:63]
  wire  _T_3884 = _T_3850 ^ _T_3882; // @[AesSbox.scala 40:63]
  wire  _T_3886 = _T_3854 ^ _T_3876; // @[AesSbox.scala 40:63]
  wire  _T_3888 = _T_3848 ^ _T_3872; // @[AesSbox.scala 40:63]
  wire  _T_3890 = matrix_3_2[7] ^ _T_3854; // @[AesSbox.scala 40:63]
  wire  _T_3892 = _T_3888 ^ _T_3856; // @[AesSbox.scala 40:63]
  wire  _T_3894 = _T_3888 ^ _T_3860; // @[AesSbox.scala 40:63]
  wire  _T_3896 = _T_3860 ^ _T_3884; // @[AesSbox.scala 40:63]
  wire  _T_3898 = _T_3878 ^ _T_3874; // @[AesSbox.scala 40:63]
  wire  _T_3900 = _T_3890 ^ _T_3880; // @[AesSbox.scala 40:63]
  wire  _T_3902 = _T_3884 & _T_3856; // @[AesSbox.scala 41:63]
  wire  _T_3904 = _T_3886 & _T_3868; // @[AesSbox.scala 41:63]
  wire  _T_3906 = _T_3870 ^ _T_3902; // @[AesSbox.scala 40:63]
  wire  _T_3908 = _T_3866 & matrix_3_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_3910 = _T_3908 ^ _T_3902; // @[AesSbox.scala 40:63]
  wire  _T_3912 = _T_3860 & _T_3888; // @[AesSbox.scala 41:63]
  wire  _T_3914 = _T_3864 & _T_3854; // @[AesSbox.scala 41:63]
  wire  _T_3916 = _T_3894 ^ _T_3912; // @[AesSbox.scala 40:63]
  wire  _T_3918 = _T_3890 & _T_3880; // @[AesSbox.scala 41:63]
  wire  _T_3920 = _T_3918 ^ _T_3912; // @[AesSbox.scala 40:63]
  wire  _T_3922 = _T_3850 & _T_3862; // @[AesSbox.scala 41:63]
  wire  _T_3924 = _T_3896 & _T_3892; // @[AesSbox.scala 41:63]
  wire  _T_3926 = _T_3924 ^ _T_3922; // @[AesSbox.scala 40:63]
  wire  _T_3928 = _T_3878 & _T_3874; // @[AesSbox.scala 41:63]
  wire  _T_3930 = _T_3928 ^ _T_3922; // @[AesSbox.scala 40:63]
  wire  _T_3932 = _T_3906 ^ _T_3904; // @[AesSbox.scala 40:63]
  wire  _T_3934 = _T_3910 ^ _T_3898; // @[AesSbox.scala 40:63]
  wire  _T_3936 = _T_3916 ^ _T_3914; // @[AesSbox.scala 40:63]
  wire  _T_3938 = _T_3920 ^ _T_3930; // @[AesSbox.scala 40:63]
  wire  _T_3940 = _T_3932 ^ _T_3926; // @[AesSbox.scala 40:63]
  wire  _T_3942 = _T_3934 ^ _T_3930; // @[AesSbox.scala 40:63]
  wire  _T_3944 = _T_3936 ^ _T_3926; // @[AesSbox.scala 40:63]
  wire  _T_3946 = _T_3938 ^ _T_3900; // @[AesSbox.scala 40:63]
  wire  _T_3948 = _T_3944 ^ _T_3946; // @[AesSbox.scala 40:63]
  wire  _T_3950 = _T_3944 & _T_3940; // @[AesSbox.scala 41:63]
  wire  _T_3952 = _T_3942 ^ _T_3950; // @[AesSbox.scala 40:63]
  wire  _T_3954 = _T_3940 ^ _T_3942; // @[AesSbox.scala 40:63]
  wire  _T_3956 = _T_3946 ^ _T_3950; // @[AesSbox.scala 40:63]
  wire  _T_3958 = _T_3956 & _T_3954; // @[AesSbox.scala 41:63]
  wire  _T_3960 = _T_3952 & _T_3948; // @[AesSbox.scala 41:63]
  wire  _T_3962 = _T_3940 & _T_3946; // @[AesSbox.scala 41:63]
  wire  _T_3964 = _T_3954 & _T_3962; // @[AesSbox.scala 41:63]
  wire  _T_3966 = _T_3954 ^ _T_3950; // @[AesSbox.scala 40:63]
  wire  _T_3968 = _T_3942 & _T_3944; // @[AesSbox.scala 41:63]
  wire  _T_3970 = _T_3948 & _T_3968; // @[AesSbox.scala 41:63]
  wire  _T_3972 = _T_3948 ^ _T_3950; // @[AesSbox.scala 40:63]
  wire  _T_3974 = _T_3942 ^ _T_3958; // @[AesSbox.scala 40:63]
  wire  _T_3976 = _T_3964 ^ _T_3966; // @[AesSbox.scala 40:63]
  wire  _T_3978 = _T_3946 ^ _T_3960; // @[AesSbox.scala 40:63]
  wire  _T_3980 = _T_3970 ^ _T_3972; // @[AesSbox.scala 40:63]
  wire  _T_3982 = _T_3976 ^ _T_3980; // @[AesSbox.scala 40:63]
  wire  _T_3984 = _T_3974 ^ _T_3978; // @[AesSbox.scala 40:63]
  wire  _T_3986 = _T_3974 ^ _T_3976; // @[AesSbox.scala 40:63]
  wire  _T_3988 = _T_3978 ^ _T_3980; // @[AesSbox.scala 40:63]
  wire  _T_3990 = _T_3984 ^ _T_3982; // @[AesSbox.scala 40:63]
  wire  _T_3992 = _T_3988 & _T_3856; // @[AesSbox.scala 41:63]
  wire  _T_3994 = _T_3980 & _T_3868; // @[AesSbox.scala 41:63]
  wire  _T_3996 = _T_3978 & matrix_3_2[0]; // @[AesSbox.scala 41:63]
  wire  _T_3998 = _T_3986 & _T_3888; // @[AesSbox.scala 41:63]
  wire  _T_4000 = _T_3976 & _T_3854; // @[AesSbox.scala 41:63]
  wire  _T_4002 = _T_3974 & _T_3880; // @[AesSbox.scala 41:63]
  wire  _T_4004 = _T_3984 & _T_3862; // @[AesSbox.scala 41:63]
  wire  _T_4006 = _T_3990 & _T_3892; // @[AesSbox.scala 41:63]
  wire  _T_4008 = _T_3982 & _T_3874; // @[AesSbox.scala 41:63]
  wire  _T_4010 = _T_3988 & _T_3884; // @[AesSbox.scala 41:63]
  wire  _T_4012 = _T_3980 & _T_3886; // @[AesSbox.scala 41:63]
  wire  _T_4014 = _T_3978 & _T_3866; // @[AesSbox.scala 41:63]
  wire  _T_4016 = _T_3986 & _T_3860; // @[AesSbox.scala 41:63]
  wire  _T_4018 = _T_3976 & _T_3864; // @[AesSbox.scala 41:63]
  wire  _T_4020 = _T_3974 & _T_3890; // @[AesSbox.scala 41:63]
  wire  _T_4022 = _T_3984 & _T_3850; // @[AesSbox.scala 41:63]
  wire  _T_4024 = _T_3990 & _T_3896; // @[AesSbox.scala 41:63]
  wire  _T_4026 = _T_3982 & _T_3878; // @[AesSbox.scala 41:63]
  wire  _T_4028 = _T_4022 ^ _T_4024; // @[AesSbox.scala 40:63]
  wire  _T_4030 = _T_4000 ^ _T_4012; // @[AesSbox.scala 40:63]
  wire  _T_4032 = _T_4006 ^ _T_4028; // @[AesSbox.scala 40:63]
  wire  _T_4034 = _T_4010 ^ _T_4030; // @[AesSbox.scala 40:63]
  wire  _T_4036 = _T_3996 ^ _T_4016; // @[AesSbox.scala 40:63]
  wire  _T_4038 = _T_3992 ^ _T_3998; // @[AesSbox.scala 40:63]
  wire  _T_4040 = _T_4028 ^ _T_4038; // @[AesSbox.scala 40:63]
  wire  _T_4042 = _T_3994 ^ _T_4034; // @[AesSbox.scala 40:63]
  wire  _T_4044 = _T_3992 ^ _T_4004; // @[AesSbox.scala 40:63]
  wire  _T_4046 = _T_4002 ^ _T_4018; // @[AesSbox.scala 40:63]
  wire  _T_4048 = _T_4008 ^ _T_4020; // @[AesSbox.scala 40:63]
  wire  _T_4050 = _T_3996 ^ _T_4042; // @[AesSbox.scala 40:63]
  wire  _T_4052 = _T_4036 ^ _T_4048; // @[AesSbox.scala 40:63]
  wire  _T_4054 = _T_4014 ^ _T_4030; // @[AesSbox.scala 40:63]
  wire  _T_4056 = _T_3998 ^ _T_4004; // @[AesSbox.scala 40:63]
  wire  _T_4058 = _T_4034 ^ _T_4056; // @[AesSbox.scala 40:63]
  wire  _T_4060 = _T_4026 ^ _T_4052; // @[AesSbox.scala 40:63]
  wire  _T_4062 = _T_4022 ^ _T_4044; // @[AesSbox.scala 40:63]
  wire  _T_4064 = _T_4036 ^ _T_4046; // @[AesSbox.scala 40:63]
  wire  _T_4065 = _T_4032 ^ _T_4058; // @[AesSbox.scala 40:63]
  wire  _T_4066 = _T_4060 ^ _T_4062; // @[AesSbox.scala 42:65]
  wire  _T_4067 = ~_T_4066; // @[AesSbox.scala 42:51]
  wire  _T_4069 = _T_4002 ^ _T_4028; // @[AesSbox.scala 40:63]
  wire  _T_4070 = _T_4040 ^ _T_4042; // @[AesSbox.scala 40:63]
  wire  _T_4071 = _T_4050 ^ _T_4069; // @[AesSbox.scala 40:63]
  wire  _T_4073 = _T_4000 ^ _T_4016; // @[AesSbox.scala 40:63]
  wire  _T_4075 = _T_4038 ^ _T_4054; // @[AesSbox.scala 40:63]
  wire  _T_4076 = _T_4040 ^ _T_4064; // @[AesSbox.scala 42:65]
  wire  _T_4077 = ~_T_4076; // @[AesSbox.scala 42:51]
  wire  _T_4079 = _T_4008 ^ _T_4046; // @[AesSbox.scala 40:63]
  wire  _T_4081 = _T_4073 ^ _T_4079; // @[AesSbox.scala 40:63]
  wire  _T_4083 = _T_4000 ^ _T_4044; // @[AesSbox.scala 40:63]
  wire  _T_4084 = _T_4032 ^ _T_4081; // @[AesSbox.scala 42:65]
  wire  _T_4085 = ~_T_4084; // @[AesSbox.scala 42:51]
  wire  _T_4087 = _T_4052 ^ _T_4075; // @[AesSbox.scala 40:63]
  wire  _T_4088 = _T_4032 ^ _T_4087; // @[AesSbox.scala 40:63]
  wire  _T_4090 = _T_4042 ^ _T_4083; // @[AesSbox.scala 40:63]
  wire  _T_4091 = _T_4032 ^ _T_4090; // @[AesSbox.scala 42:65]
  wire  _T_4092 = ~_T_4091; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_1_2 = {_T_4065,_T_4092,_T_4067,_T_4070,_T_4071,_T_4088,_T_4085,_T_4077}; // @[Cat.scala 29:58]
  wire  _T_4117 = matrix_3_3[1] ^ matrix_3_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_4119 = matrix_3_3[4] ^ matrix_3_3[7]; // @[AesSbox.scala 40:63]
  wire  _T_4121 = matrix_3_3[6] ^ matrix_3_3[5]; // @[AesSbox.scala 40:63]
  wire  _T_4123 = matrix_3_3[0] ^ _T_4121; // @[AesSbox.scala 40:63]
  wire  _T_4125 = _T_4117 ^ _T_4119; // @[AesSbox.scala 40:63]
  wire  _T_4127 = matrix_3_3[6] ^ matrix_3_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_4129 = matrix_3_3[7] ^ matrix_3_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_4131 = _T_4117 ^ _T_4127; // @[AesSbox.scala 40:63]
  wire  _T_4133 = matrix_3_3[1] ^ _T_4123; // @[AesSbox.scala 40:63]
  wire  _T_4135 = matrix_3_3[4] ^ _T_4123; // @[AesSbox.scala 40:63]
  wire  _T_4137 = matrix_3_3[0] ^ _T_4125; // @[AesSbox.scala 40:63]
  wire  _T_4139 = _T_4125 ^ _T_4127; // @[AesSbox.scala 40:63]
  wire  _T_4141 = matrix_3_3[5] ^ matrix_3_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_4143 = _T_4121 ^ _T_4125; // @[AesSbox.scala 40:63]
  wire  _T_4145 = matrix_3_3[2] ^ _T_4129; // @[AesSbox.scala 40:63]
  wire  _T_4147 = matrix_3_3[7] ^ matrix_3_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_4149 = matrix_3_3[0] ^ _T_4131; // @[AesSbox.scala 40:63]
  wire  _T_4151 = matrix_3_3[1] ^ matrix_3_3[2]; // @[AesSbox.scala 40:63]
  wire  _T_4153 = _T_4119 ^ _T_4151; // @[AesSbox.scala 40:63]
  wire  _T_4155 = _T_4123 ^ _T_4145; // @[AesSbox.scala 40:63]
  wire  _T_4157 = _T_4117 ^ _T_4141; // @[AesSbox.scala 40:63]
  wire  _T_4159 = matrix_3_3[7] ^ _T_4123; // @[AesSbox.scala 40:63]
  wire  _T_4161 = _T_4157 ^ _T_4125; // @[AesSbox.scala 40:63]
  wire  _T_4163 = _T_4157 ^ _T_4129; // @[AesSbox.scala 40:63]
  wire  _T_4165 = _T_4129 ^ _T_4153; // @[AesSbox.scala 40:63]
  wire  _T_4167 = _T_4147 ^ _T_4143; // @[AesSbox.scala 40:63]
  wire  _T_4169 = _T_4159 ^ _T_4149; // @[AesSbox.scala 40:63]
  wire  _T_4171 = _T_4153 & _T_4125; // @[AesSbox.scala 41:63]
  wire  _T_4173 = _T_4155 & _T_4137; // @[AesSbox.scala 41:63]
  wire  _T_4175 = _T_4139 ^ _T_4171; // @[AesSbox.scala 40:63]
  wire  _T_4177 = _T_4135 & matrix_3_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_4179 = _T_4177 ^ _T_4171; // @[AesSbox.scala 40:63]
  wire  _T_4181 = _T_4129 & _T_4157; // @[AesSbox.scala 41:63]
  wire  _T_4183 = _T_4133 & _T_4123; // @[AesSbox.scala 41:63]
  wire  _T_4185 = _T_4163 ^ _T_4181; // @[AesSbox.scala 40:63]
  wire  _T_4187 = _T_4159 & _T_4149; // @[AesSbox.scala 41:63]
  wire  _T_4189 = _T_4187 ^ _T_4181; // @[AesSbox.scala 40:63]
  wire  _T_4191 = _T_4119 & _T_4131; // @[AesSbox.scala 41:63]
  wire  _T_4193 = _T_4165 & _T_4161; // @[AesSbox.scala 41:63]
  wire  _T_4195 = _T_4193 ^ _T_4191; // @[AesSbox.scala 40:63]
  wire  _T_4197 = _T_4147 & _T_4143; // @[AesSbox.scala 41:63]
  wire  _T_4199 = _T_4197 ^ _T_4191; // @[AesSbox.scala 40:63]
  wire  _T_4201 = _T_4175 ^ _T_4173; // @[AesSbox.scala 40:63]
  wire  _T_4203 = _T_4179 ^ _T_4167; // @[AesSbox.scala 40:63]
  wire  _T_4205 = _T_4185 ^ _T_4183; // @[AesSbox.scala 40:63]
  wire  _T_4207 = _T_4189 ^ _T_4199; // @[AesSbox.scala 40:63]
  wire  _T_4209 = _T_4201 ^ _T_4195; // @[AesSbox.scala 40:63]
  wire  _T_4211 = _T_4203 ^ _T_4199; // @[AesSbox.scala 40:63]
  wire  _T_4213 = _T_4205 ^ _T_4195; // @[AesSbox.scala 40:63]
  wire  _T_4215 = _T_4207 ^ _T_4169; // @[AesSbox.scala 40:63]
  wire  _T_4217 = _T_4213 ^ _T_4215; // @[AesSbox.scala 40:63]
  wire  _T_4219 = _T_4213 & _T_4209; // @[AesSbox.scala 41:63]
  wire  _T_4221 = _T_4211 ^ _T_4219; // @[AesSbox.scala 40:63]
  wire  _T_4223 = _T_4209 ^ _T_4211; // @[AesSbox.scala 40:63]
  wire  _T_4225 = _T_4215 ^ _T_4219; // @[AesSbox.scala 40:63]
  wire  _T_4227 = _T_4225 & _T_4223; // @[AesSbox.scala 41:63]
  wire  _T_4229 = _T_4221 & _T_4217; // @[AesSbox.scala 41:63]
  wire  _T_4231 = _T_4209 & _T_4215; // @[AesSbox.scala 41:63]
  wire  _T_4233 = _T_4223 & _T_4231; // @[AesSbox.scala 41:63]
  wire  _T_4235 = _T_4223 ^ _T_4219; // @[AesSbox.scala 40:63]
  wire  _T_4237 = _T_4211 & _T_4213; // @[AesSbox.scala 41:63]
  wire  _T_4239 = _T_4217 & _T_4237; // @[AesSbox.scala 41:63]
  wire  _T_4241 = _T_4217 ^ _T_4219; // @[AesSbox.scala 40:63]
  wire  _T_4243 = _T_4211 ^ _T_4227; // @[AesSbox.scala 40:63]
  wire  _T_4245 = _T_4233 ^ _T_4235; // @[AesSbox.scala 40:63]
  wire  _T_4247 = _T_4215 ^ _T_4229; // @[AesSbox.scala 40:63]
  wire  _T_4249 = _T_4239 ^ _T_4241; // @[AesSbox.scala 40:63]
  wire  _T_4251 = _T_4245 ^ _T_4249; // @[AesSbox.scala 40:63]
  wire  _T_4253 = _T_4243 ^ _T_4247; // @[AesSbox.scala 40:63]
  wire  _T_4255 = _T_4243 ^ _T_4245; // @[AesSbox.scala 40:63]
  wire  _T_4257 = _T_4247 ^ _T_4249; // @[AesSbox.scala 40:63]
  wire  _T_4259 = _T_4253 ^ _T_4251; // @[AesSbox.scala 40:63]
  wire  _T_4261 = _T_4257 & _T_4125; // @[AesSbox.scala 41:63]
  wire  _T_4263 = _T_4249 & _T_4137; // @[AesSbox.scala 41:63]
  wire  _T_4265 = _T_4247 & matrix_3_3[0]; // @[AesSbox.scala 41:63]
  wire  _T_4267 = _T_4255 & _T_4157; // @[AesSbox.scala 41:63]
  wire  _T_4269 = _T_4245 & _T_4123; // @[AesSbox.scala 41:63]
  wire  _T_4271 = _T_4243 & _T_4149; // @[AesSbox.scala 41:63]
  wire  _T_4273 = _T_4253 & _T_4131; // @[AesSbox.scala 41:63]
  wire  _T_4275 = _T_4259 & _T_4161; // @[AesSbox.scala 41:63]
  wire  _T_4277 = _T_4251 & _T_4143; // @[AesSbox.scala 41:63]
  wire  _T_4279 = _T_4257 & _T_4153; // @[AesSbox.scala 41:63]
  wire  _T_4281 = _T_4249 & _T_4155; // @[AesSbox.scala 41:63]
  wire  _T_4283 = _T_4247 & _T_4135; // @[AesSbox.scala 41:63]
  wire  _T_4285 = _T_4255 & _T_4129; // @[AesSbox.scala 41:63]
  wire  _T_4287 = _T_4245 & _T_4133; // @[AesSbox.scala 41:63]
  wire  _T_4289 = _T_4243 & _T_4159; // @[AesSbox.scala 41:63]
  wire  _T_4291 = _T_4253 & _T_4119; // @[AesSbox.scala 41:63]
  wire  _T_4293 = _T_4259 & _T_4165; // @[AesSbox.scala 41:63]
  wire  _T_4295 = _T_4251 & _T_4147; // @[AesSbox.scala 41:63]
  wire  _T_4297 = _T_4291 ^ _T_4293; // @[AesSbox.scala 40:63]
  wire  _T_4299 = _T_4269 ^ _T_4281; // @[AesSbox.scala 40:63]
  wire  _T_4301 = _T_4275 ^ _T_4297; // @[AesSbox.scala 40:63]
  wire  _T_4303 = _T_4279 ^ _T_4299; // @[AesSbox.scala 40:63]
  wire  _T_4305 = _T_4265 ^ _T_4285; // @[AesSbox.scala 40:63]
  wire  _T_4307 = _T_4261 ^ _T_4267; // @[AesSbox.scala 40:63]
  wire  _T_4309 = _T_4297 ^ _T_4307; // @[AesSbox.scala 40:63]
  wire  _T_4311 = _T_4263 ^ _T_4303; // @[AesSbox.scala 40:63]
  wire  _T_4313 = _T_4261 ^ _T_4273; // @[AesSbox.scala 40:63]
  wire  _T_4315 = _T_4271 ^ _T_4287; // @[AesSbox.scala 40:63]
  wire  _T_4317 = _T_4277 ^ _T_4289; // @[AesSbox.scala 40:63]
  wire  _T_4319 = _T_4265 ^ _T_4311; // @[AesSbox.scala 40:63]
  wire  _T_4321 = _T_4305 ^ _T_4317; // @[AesSbox.scala 40:63]
  wire  _T_4323 = _T_4283 ^ _T_4299; // @[AesSbox.scala 40:63]
  wire  _T_4325 = _T_4267 ^ _T_4273; // @[AesSbox.scala 40:63]
  wire  _T_4327 = _T_4303 ^ _T_4325; // @[AesSbox.scala 40:63]
  wire  _T_4329 = _T_4295 ^ _T_4321; // @[AesSbox.scala 40:63]
  wire  _T_4331 = _T_4291 ^ _T_4313; // @[AesSbox.scala 40:63]
  wire  _T_4333 = _T_4305 ^ _T_4315; // @[AesSbox.scala 40:63]
  wire  _T_4334 = _T_4301 ^ _T_4327; // @[AesSbox.scala 40:63]
  wire  _T_4335 = _T_4329 ^ _T_4331; // @[AesSbox.scala 42:65]
  wire  _T_4336 = ~_T_4335; // @[AesSbox.scala 42:51]
  wire  _T_4338 = _T_4271 ^ _T_4297; // @[AesSbox.scala 40:63]
  wire  _T_4339 = _T_4309 ^ _T_4311; // @[AesSbox.scala 40:63]
  wire  _T_4340 = _T_4319 ^ _T_4338; // @[AesSbox.scala 40:63]
  wire  _T_4342 = _T_4269 ^ _T_4285; // @[AesSbox.scala 40:63]
  wire  _T_4344 = _T_4307 ^ _T_4323; // @[AesSbox.scala 40:63]
  wire  _T_4345 = _T_4309 ^ _T_4333; // @[AesSbox.scala 42:65]
  wire  _T_4346 = ~_T_4345; // @[AesSbox.scala 42:51]
  wire  _T_4348 = _T_4277 ^ _T_4315; // @[AesSbox.scala 40:63]
  wire  _T_4350 = _T_4342 ^ _T_4348; // @[AesSbox.scala 40:63]
  wire  _T_4352 = _T_4269 ^ _T_4313; // @[AesSbox.scala 40:63]
  wire  _T_4353 = _T_4301 ^ _T_4350; // @[AesSbox.scala 42:65]
  wire  _T_4354 = ~_T_4353; // @[AesSbox.scala 42:51]
  wire  _T_4356 = _T_4321 ^ _T_4344; // @[AesSbox.scala 40:63]
  wire  _T_4357 = _T_4301 ^ _T_4356; // @[AesSbox.scala 40:63]
  wire  _T_4359 = _T_4311 ^ _T_4352; // @[AesSbox.scala 40:63]
  wire  _T_4360 = _T_4301 ^ _T_4359; // @[AesSbox.scala 42:65]
  wire  _T_4361 = ~_T_4360; // @[AesSbox.scala 42:51]
  wire [7:0] roundPart1_0_3 = {_T_4334,_T_4361,_T_4336,_T_4339,_T_4340,_T_4357,_T_4354,_T_4346}; // @[Cat.scala 29:58]
  wire [7:0] roundPart2_0_0 = MixColsModule_io_out_0_0 ^ io_keys_0_0_0; // @[AesComponents.scala 57:30]
  wire [7:0] roundPart2_0_1 = MixColsModule_io_out_0_1 ^ io_keys_0_0_1; // @[AesComponents.scala 57:51]
  wire [7:0] roundPart2_0_2 = MixColsModule_io_out_0_2 ^ io_keys_0_0_2; // @[AesComponents.scala 57:72]
  wire [7:0] roundPart2_0_3 = MixColsModule_io_out_0_3 ^ io_keys_0_0_3; // @[AesComponents.scala 57:93]
  wire [7:0] roundPart2_1_0 = MixColsModule_io_out_1_0 ^ io_keys_0_1_0; // @[AesComponents.scala 58:30]
  wire [7:0] roundPart2_1_1 = MixColsModule_io_out_1_1 ^ io_keys_0_1_1; // @[AesComponents.scala 58:51]
  wire [7:0] roundPart2_1_2 = MixColsModule_io_out_1_2 ^ io_keys_0_1_2; // @[AesComponents.scala 58:72]
  wire [7:0] roundPart2_1_3 = MixColsModule_io_out_1_3 ^ io_keys_0_1_3; // @[AesComponents.scala 58:93]
  wire [7:0] roundPart2_2_0 = MixColsModule_io_out_2_0 ^ io_keys_0_2_0; // @[AesComponents.scala 59:30]
  wire [7:0] roundPart2_2_1 = MixColsModule_io_out_2_1 ^ io_keys_0_2_1; // @[AesComponents.scala 59:51]
  wire [7:0] roundPart2_2_2 = MixColsModule_io_out_2_2 ^ io_keys_0_2_2; // @[AesComponents.scala 59:72]
  wire [7:0] roundPart2_2_3 = MixColsModule_io_out_2_3 ^ io_keys_0_2_3; // @[AesComponents.scala 59:93]
  wire [7:0] roundPart2_3_0 = MixColsModule_io_out_3_0 ^ io_keys_0_3_0; // @[AesComponents.scala 60:30]
  wire [7:0] roundPart2_3_1 = MixColsModule_io_out_3_1 ^ io_keys_0_3_1; // @[AesComponents.scala 60:51]
  wire [7:0] roundPart2_3_2 = MixColsModule_io_out_3_2 ^ io_keys_0_3_2; // @[AesComponents.scala 60:72]
  wire [7:0] roundPart2_3_3 = MixColsModule_io_out_3_3 ^ io_keys_0_3_3; // @[AesComponents.scala 60:93]
  wire [7:0] roundPart2_last_0_0 = matrix_0_0 ^ io_keys_0_0_0; // @[AesComponents.scala 57:30]
  wire [7:0] roundPart2_last_0_1 = matrix_0_1 ^ io_keys_0_0_1; // @[AesComponents.scala 57:51]
  wire [7:0] roundPart2_last_0_2 = matrix_0_2 ^ io_keys_0_0_2; // @[AesComponents.scala 57:72]
  wire [7:0] roundPart2_last_0_3 = matrix_0_3 ^ io_keys_0_0_3; // @[AesComponents.scala 57:93]
  wire [7:0] roundPart2_last_1_0 = matrix_1_0 ^ io_keys_0_1_0; // @[AesComponents.scala 58:30]
  wire [7:0] roundPart2_last_1_1 = matrix_1_1 ^ io_keys_0_1_1; // @[AesComponents.scala 58:51]
  wire [7:0] roundPart2_last_1_2 = matrix_1_2 ^ io_keys_0_1_2; // @[AesComponents.scala 58:72]
  wire [7:0] roundPart2_last_1_3 = matrix_1_3 ^ io_keys_0_1_3; // @[AesComponents.scala 58:93]
  wire [7:0] roundPart2_last_2_0 = matrix_2_0 ^ io_keys_0_2_0; // @[AesComponents.scala 59:30]
  wire [7:0] roundPart2_last_2_1 = matrix_2_1 ^ io_keys_0_2_1; // @[AesComponents.scala 59:51]
  wire [7:0] roundPart2_last_2_2 = matrix_2_2 ^ io_keys_0_2_2; // @[AesComponents.scala 59:72]
  wire [7:0] roundPart2_last_2_3 = matrix_2_3 ^ io_keys_0_2_3; // @[AesComponents.scala 59:93]
  wire [7:0] roundPart2_last_3_0 = matrix_3_0 ^ io_keys_0_3_0; // @[AesComponents.scala 60:30]
  wire [7:0] roundPart2_last_3_1 = matrix_3_1 ^ io_keys_0_3_1; // @[AesComponents.scala 60:51]
  wire [7:0] roundPart2_last_3_2 = matrix_3_2 ^ io_keys_0_3_2; // @[AesComponents.scala 60:72]
  wire [7:0] roundPart2_last_3_3 = matrix_3_3 ^ io_keys_0_3_3; // @[AesComponents.scala 60:93]
  wire  _T_4415 = io_ready & io_dataValid; // @[AesEncrypt.scala 75:20]
  wire  _T_4417 = state == 6'h1d; // @[AesEncrypt.scala 82:41]
  wire  _T_4418 = state == 6'h15; // @[AesEncrypt.scala 82:57]
  wire  _T_4419 = io_aes256 ? _T_4417 : _T_4418; // @[AesEncrypt.scala 82:23]
  wire  _T_4421 = ~state[0]; // @[AesEncrypt.scala 84:24]
  wire  _GEN_34 = _T_4421 ? _T_4415 : 1'h1; // @[AesEncrypt.scala 84:33]
  wire [5:0] _T_4424 = state + 6'h1; // @[AesEncrypt.scala 91:24]
  MixColsModule MixColsModule ( // @[AesComponents.scala 91:35]
    .io_in_0_0(MixColsModule_io_in_0_0),
    .io_in_0_1(MixColsModule_io_in_0_1),
    .io_in_0_2(MixColsModule_io_in_0_2),
    .io_in_0_3(MixColsModule_io_in_0_3),
    .io_in_1_0(MixColsModule_io_in_1_0),
    .io_in_1_1(MixColsModule_io_in_1_1),
    .io_in_1_2(MixColsModule_io_in_1_2),
    .io_in_1_3(MixColsModule_io_in_1_3),
    .io_in_2_0(MixColsModule_io_in_2_0),
    .io_in_2_1(MixColsModule_io_in_2_1),
    .io_in_2_2(MixColsModule_io_in_2_2),
    .io_in_2_3(MixColsModule_io_in_2_3),
    .io_in_3_0(MixColsModule_io_in_3_0),
    .io_in_3_1(MixColsModule_io_in_3_1),
    .io_in_3_2(MixColsModule_io_in_3_2),
    .io_in_3_3(MixColsModule_io_in_3_3),
    .io_out_0_0(MixColsModule_io_out_0_0),
    .io_out_0_1(MixColsModule_io_out_0_1),
    .io_out_0_2(MixColsModule_io_out_0_2),
    .io_out_0_3(MixColsModule_io_out_0_3),
    .io_out_1_0(MixColsModule_io_out_1_0),
    .io_out_1_1(MixColsModule_io_out_1_1),
    .io_out_1_2(MixColsModule_io_out_1_2),
    .io_out_1_3(MixColsModule_io_out_1_3),
    .io_out_2_0(MixColsModule_io_out_2_0),
    .io_out_2_1(MixColsModule_io_out_2_1),
    .io_out_2_2(MixColsModule_io_out_2_2),
    .io_out_2_3(MixColsModule_io_out_2_3),
    .io_out_3_0(MixColsModule_io_out_3_0),
    .io_out_3_1(MixColsModule_io_out_3_1),
    .io_out_3_2(MixColsModule_io_out_3_2),
    .io_out_3_3(MixColsModule_io_out_3_3)
  );
  assign io_shiftCyc = _T_6 | io_dataValid; // @[AesEncrypt.scala 60:17]
  assign io_shift = _T_6 ? _GEN_34 : _T_4415; // @[AesEncrypt.scala 61:14 AesEncrypt.scala 78:18 AesEncrypt.scala 88:22]
  assign io_ready = _T_2 | _T_3; // @[AesEncrypt.scala 56:14]
  assign io_dataOut = {_T_23,_T_16}; // @[AesEncrypt.scala 65:16]
  assign io_ivOut = io_dataOut; // @[AesEncrypt.scala 66:14]
  assign io_outputValid = state == 6'h1e; // @[AesEncrypt.scala 57:20]
  assign MixColsModule_io_in_0_0 = matrix_0_0; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_0_1 = matrix_0_1; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_0_2 = matrix_0_2; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_0_3 = matrix_0_3; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_0 = matrix_1_0; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_1 = matrix_1_1; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_2 = matrix_1_2; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_3 = matrix_1_3; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_0 = matrix_2_0; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_1 = matrix_2_1; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_2 = matrix_2_2; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_3 = matrix_2_3; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_0 = matrix_3_0; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_1 = matrix_3_1; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_2 = matrix_3_2; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_3 = matrix_3_3; // @[AesComponents.scala 92:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  matrix_0_0 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  matrix_0_1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  matrix_0_2 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  matrix_0_3 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  matrix_1_0 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  matrix_1_1 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  matrix_1_2 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  matrix_1_3 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  matrix_2_0 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  matrix_2_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  matrix_2_2 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  matrix_2_3 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  matrix_3_0 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  matrix_3_1 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  matrix_3_2 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  matrix_3_3 = _RAND_16[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 6'h1;
    end else if (_T_6) begin
      if (_T_4419) begin
        state <= 6'h1e;
      end else begin
        state <= _T_4424;
      end
    end else if (_T_4415) begin
      state <= 6'h2;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_0_0 <= roundPart1_0_0;
      end else if (_T_4419) begin
        matrix_0_0 <= roundPart2_last_0_0;
      end else begin
        matrix_0_0 <= roundPart2_0_0;
      end
    end else if (_T_4415) begin
      matrix_0_0 <= initOut_0_0;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_0_1 <= roundPart1_0_1;
      end else if (_T_4419) begin
        matrix_0_1 <= roundPart2_last_0_1;
      end else begin
        matrix_0_1 <= roundPart2_0_1;
      end
    end else if (_T_4415) begin
      matrix_0_1 <= initOut_0_1;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_0_2 <= roundPart1_0_2;
      end else if (_T_4419) begin
        matrix_0_2 <= roundPart2_last_0_2;
      end else begin
        matrix_0_2 <= roundPart2_0_2;
      end
    end else if (_T_4415) begin
      matrix_0_2 <= initOut_0_2;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_0_3 <= roundPart1_0_3;
      end else if (_T_4419) begin
        matrix_0_3 <= roundPart2_last_0_3;
      end else begin
        matrix_0_3 <= roundPart2_0_3;
      end
    end else if (_T_4415) begin
      matrix_0_3 <= initOut_0_3;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_1_0 <= roundPart1_1_0;
      end else if (_T_4419) begin
        matrix_1_0 <= roundPart2_last_1_0;
      end else begin
        matrix_1_0 <= roundPart2_1_0;
      end
    end else if (_T_4415) begin
      matrix_1_0 <= initOut_1_0;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_1_1 <= roundPart1_1_1;
      end else if (_T_4419) begin
        matrix_1_1 <= roundPart2_last_1_1;
      end else begin
        matrix_1_1 <= roundPart2_1_1;
      end
    end else if (_T_4415) begin
      matrix_1_1 <= initOut_1_1;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_1_2 <= roundPart1_1_2;
      end else if (_T_4419) begin
        matrix_1_2 <= roundPart2_last_1_2;
      end else begin
        matrix_1_2 <= roundPart2_1_2;
      end
    end else if (_T_4415) begin
      matrix_1_2 <= initOut_1_2;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_1_3 <= roundPart1_1_3;
      end else if (_T_4419) begin
        matrix_1_3 <= roundPart2_last_1_3;
      end else begin
        matrix_1_3 <= roundPart2_1_3;
      end
    end else if (_T_4415) begin
      matrix_1_3 <= initOut_1_3;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_2_0 <= roundPart1_2_0;
      end else if (_T_4419) begin
        matrix_2_0 <= roundPart2_last_2_0;
      end else begin
        matrix_2_0 <= roundPart2_2_0;
      end
    end else if (_T_4415) begin
      matrix_2_0 <= initOut_2_0;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_2_1 <= roundPart1_2_1;
      end else if (_T_4419) begin
        matrix_2_1 <= roundPart2_last_2_1;
      end else begin
        matrix_2_1 <= roundPart2_2_1;
      end
    end else if (_T_4415) begin
      matrix_2_1 <= initOut_2_1;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_2_2 <= roundPart1_2_2;
      end else if (_T_4419) begin
        matrix_2_2 <= roundPart2_last_2_2;
      end else begin
        matrix_2_2 <= roundPart2_2_2;
      end
    end else if (_T_4415) begin
      matrix_2_2 <= initOut_2_2;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_2_3 <= roundPart1_2_3;
      end else if (_T_4419) begin
        matrix_2_3 <= roundPart2_last_2_3;
      end else begin
        matrix_2_3 <= roundPart2_2_3;
      end
    end else if (_T_4415) begin
      matrix_2_3 <= initOut_2_3;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_3_0 <= roundPart1_3_0;
      end else if (_T_4419) begin
        matrix_3_0 <= roundPart2_last_3_0;
      end else begin
        matrix_3_0 <= roundPart2_3_0;
      end
    end else if (_T_4415) begin
      matrix_3_0 <= initOut_3_0;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_3_1 <= roundPart1_3_1;
      end else if (_T_4419) begin
        matrix_3_1 <= roundPart2_last_3_1;
      end else begin
        matrix_3_1 <= roundPart2_3_1;
      end
    end else if (_T_4415) begin
      matrix_3_1 <= initOut_3_1;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_3_2 <= roundPart1_3_2;
      end else if (_T_4419) begin
        matrix_3_2 <= roundPart2_last_3_2;
      end else begin
        matrix_3_2 <= roundPart2_3_2;
      end
    end else if (_T_4415) begin
      matrix_3_2 <= initOut_3_2;
    end
    if (_T_6) begin
      if (_T_4421) begin
        matrix_3_3 <= roundPart1_3_3;
      end else if (_T_4419) begin
        matrix_3_3 <= roundPart2_last_3_3;
      end else begin
        matrix_3_3 <= roundPart2_3_3;
      end
    end else if (_T_4415) begin
      matrix_3_3 <= initOut_3_3;
    end
  end
endmodule
module AesDecrypt(
  input          clock,
  input          reset,
  input  [127:0] io_dataIn,
  input  [127:0] io_ivIn,
  input          io_dataValid,
  input  [7:0]   io_keys_0_0_0,
  input  [7:0]   io_keys_0_0_1,
  input  [7:0]   io_keys_0_0_2,
  input  [7:0]   io_keys_0_0_3,
  input  [7:0]   io_keys_0_1_0,
  input  [7:0]   io_keys_0_1_1,
  input  [7:0]   io_keys_0_1_2,
  input  [7:0]   io_keys_0_1_3,
  input  [7:0]   io_keys_0_2_0,
  input  [7:0]   io_keys_0_2_1,
  input  [7:0]   io_keys_0_2_2,
  input  [7:0]   io_keys_0_2_3,
  input  [7:0]   io_keys_0_3_0,
  input  [7:0]   io_keys_0_3_1,
  input  [7:0]   io_keys_0_3_2,
  input  [7:0]   io_keys_0_3_3,
  input  [7:0]   io_keys_1_0_0,
  input  [7:0]   io_keys_1_0_1,
  input  [7:0]   io_keys_1_0_2,
  input  [7:0]   io_keys_1_0_3,
  input  [7:0]   io_keys_1_1_0,
  input  [7:0]   io_keys_1_1_1,
  input  [7:0]   io_keys_1_1_2,
  input  [7:0]   io_keys_1_1_3,
  input  [7:0]   io_keys_1_2_0,
  input  [7:0]   io_keys_1_2_1,
  input  [7:0]   io_keys_1_2_2,
  input  [7:0]   io_keys_1_2_3,
  input  [7:0]   io_keys_1_3_0,
  input  [7:0]   io_keys_1_3_1,
  input  [7:0]   io_keys_1_3_2,
  input  [7:0]   io_keys_1_3_3,
  input  [7:0]   io_keys_2_0_0,
  input  [7:0]   io_keys_2_0_1,
  input  [7:0]   io_keys_2_0_2,
  input  [7:0]   io_keys_2_0_3,
  input  [7:0]   io_keys_2_1_0,
  input  [7:0]   io_keys_2_1_1,
  input  [7:0]   io_keys_2_1_2,
  input  [7:0]   io_keys_2_1_3,
  input  [7:0]   io_keys_2_2_0,
  input  [7:0]   io_keys_2_2_1,
  input  [7:0]   io_keys_2_2_2,
  input  [7:0]   io_keys_2_2_3,
  input  [7:0]   io_keys_2_3_0,
  input  [7:0]   io_keys_2_3_1,
  input  [7:0]   io_keys_2_3_2,
  input  [7:0]   io_keys_2_3_3,
  input  [7:0]   io_keys_3_0_0,
  input  [7:0]   io_keys_3_0_1,
  input  [7:0]   io_keys_3_0_2,
  input  [7:0]   io_keys_3_0_3,
  input  [7:0]   io_keys_3_1_0,
  input  [7:0]   io_keys_3_1_1,
  input  [7:0]   io_keys_3_1_2,
  input  [7:0]   io_keys_3_1_3,
  input  [7:0]   io_keys_3_2_0,
  input  [7:0]   io_keys_3_2_1,
  input  [7:0]   io_keys_3_2_2,
  input  [7:0]   io_keys_3_2_3,
  input  [7:0]   io_keys_3_3_0,
  input  [7:0]   io_keys_3_3_1,
  input  [7:0]   io_keys_3_3_2,
  input  [7:0]   io_keys_3_3_3,
  input  [7:0]   io_keys_4_0_0,
  input  [7:0]   io_keys_4_0_1,
  input  [7:0]   io_keys_4_0_2,
  input  [7:0]   io_keys_4_0_3,
  input  [7:0]   io_keys_4_1_0,
  input  [7:0]   io_keys_4_1_1,
  input  [7:0]   io_keys_4_1_2,
  input  [7:0]   io_keys_4_1_3,
  input  [7:0]   io_keys_4_2_0,
  input  [7:0]   io_keys_4_2_1,
  input  [7:0]   io_keys_4_2_2,
  input  [7:0]   io_keys_4_2_3,
  input  [7:0]   io_keys_4_3_0,
  input  [7:0]   io_keys_4_3_1,
  input  [7:0]   io_keys_4_3_2,
  input  [7:0]   io_keys_4_3_3,
  input  [7:0]   io_keys_5_0_0,
  input  [7:0]   io_keys_5_0_1,
  input  [7:0]   io_keys_5_0_2,
  input  [7:0]   io_keys_5_0_3,
  input  [7:0]   io_keys_5_1_0,
  input  [7:0]   io_keys_5_1_1,
  input  [7:0]   io_keys_5_1_2,
  input  [7:0]   io_keys_5_1_3,
  input  [7:0]   io_keys_5_2_0,
  input  [7:0]   io_keys_5_2_1,
  input  [7:0]   io_keys_5_2_2,
  input  [7:0]   io_keys_5_2_3,
  input  [7:0]   io_keys_5_3_0,
  input  [7:0]   io_keys_5_3_1,
  input  [7:0]   io_keys_5_3_2,
  input  [7:0]   io_keys_5_3_3,
  input  [7:0]   io_keys_6_0_0,
  input  [7:0]   io_keys_6_0_1,
  input  [7:0]   io_keys_6_0_2,
  input  [7:0]   io_keys_6_0_3,
  input  [7:0]   io_keys_6_1_0,
  input  [7:0]   io_keys_6_1_1,
  input  [7:0]   io_keys_6_1_2,
  input  [7:0]   io_keys_6_1_3,
  input  [7:0]   io_keys_6_2_0,
  input  [7:0]   io_keys_6_2_1,
  input  [7:0]   io_keys_6_2_2,
  input  [7:0]   io_keys_6_2_3,
  input  [7:0]   io_keys_6_3_0,
  input  [7:0]   io_keys_6_3_1,
  input  [7:0]   io_keys_6_3_2,
  input  [7:0]   io_keys_6_3_3,
  input  [7:0]   io_keys_7_0_0,
  input  [7:0]   io_keys_7_0_1,
  input  [7:0]   io_keys_7_0_2,
  input  [7:0]   io_keys_7_0_3,
  input  [7:0]   io_keys_7_1_0,
  input  [7:0]   io_keys_7_1_1,
  input  [7:0]   io_keys_7_1_2,
  input  [7:0]   io_keys_7_1_3,
  input  [7:0]   io_keys_7_2_0,
  input  [7:0]   io_keys_7_2_1,
  input  [7:0]   io_keys_7_2_2,
  input  [7:0]   io_keys_7_2_3,
  input  [7:0]   io_keys_7_3_0,
  input  [7:0]   io_keys_7_3_1,
  input  [7:0]   io_keys_7_3_2,
  input  [7:0]   io_keys_7_3_3,
  input  [7:0]   io_keys_8_0_0,
  input  [7:0]   io_keys_8_0_1,
  input  [7:0]   io_keys_8_0_2,
  input  [7:0]   io_keys_8_0_3,
  input  [7:0]   io_keys_8_1_0,
  input  [7:0]   io_keys_8_1_1,
  input  [7:0]   io_keys_8_1_2,
  input  [7:0]   io_keys_8_1_3,
  input  [7:0]   io_keys_8_2_0,
  input  [7:0]   io_keys_8_2_1,
  input  [7:0]   io_keys_8_2_2,
  input  [7:0]   io_keys_8_2_3,
  input  [7:0]   io_keys_8_3_0,
  input  [7:0]   io_keys_8_3_1,
  input  [7:0]   io_keys_8_3_2,
  input  [7:0]   io_keys_8_3_3,
  input  [7:0]   io_keys_9_0_0,
  input  [7:0]   io_keys_9_0_1,
  input  [7:0]   io_keys_9_0_2,
  input  [7:0]   io_keys_9_0_3,
  input  [7:0]   io_keys_9_1_0,
  input  [7:0]   io_keys_9_1_1,
  input  [7:0]   io_keys_9_1_2,
  input  [7:0]   io_keys_9_1_3,
  input  [7:0]   io_keys_9_2_0,
  input  [7:0]   io_keys_9_2_1,
  input  [7:0]   io_keys_9_2_2,
  input  [7:0]   io_keys_9_2_3,
  input  [7:0]   io_keys_9_3_0,
  input  [7:0]   io_keys_9_3_1,
  input  [7:0]   io_keys_9_3_2,
  input  [7:0]   io_keys_9_3_3,
  input  [7:0]   io_keys_10_0_0,
  input  [7:0]   io_keys_10_0_1,
  input  [7:0]   io_keys_10_0_2,
  input  [7:0]   io_keys_10_0_3,
  input  [7:0]   io_keys_10_1_0,
  input  [7:0]   io_keys_10_1_1,
  input  [7:0]   io_keys_10_1_2,
  input  [7:0]   io_keys_10_1_3,
  input  [7:0]   io_keys_10_2_0,
  input  [7:0]   io_keys_10_2_1,
  input  [7:0]   io_keys_10_2_2,
  input  [7:0]   io_keys_10_2_3,
  input  [7:0]   io_keys_10_3_0,
  input  [7:0]   io_keys_10_3_1,
  input  [7:0]   io_keys_10_3_2,
  input  [7:0]   io_keys_10_3_3,
  input  [7:0]   io_keys_11_0_0,
  input  [7:0]   io_keys_11_0_1,
  input  [7:0]   io_keys_11_0_2,
  input  [7:0]   io_keys_11_0_3,
  input  [7:0]   io_keys_11_1_0,
  input  [7:0]   io_keys_11_1_1,
  input  [7:0]   io_keys_11_1_2,
  input  [7:0]   io_keys_11_1_3,
  input  [7:0]   io_keys_11_2_0,
  input  [7:0]   io_keys_11_2_1,
  input  [7:0]   io_keys_11_2_2,
  input  [7:0]   io_keys_11_2_3,
  input  [7:0]   io_keys_11_3_0,
  input  [7:0]   io_keys_11_3_1,
  input  [7:0]   io_keys_11_3_2,
  input  [7:0]   io_keys_11_3_3,
  input  [7:0]   io_keys_12_0_0,
  input  [7:0]   io_keys_12_0_1,
  input  [7:0]   io_keys_12_0_2,
  input  [7:0]   io_keys_12_0_3,
  input  [7:0]   io_keys_12_1_0,
  input  [7:0]   io_keys_12_1_1,
  input  [7:0]   io_keys_12_1_2,
  input  [7:0]   io_keys_12_1_3,
  input  [7:0]   io_keys_12_2_0,
  input  [7:0]   io_keys_12_2_1,
  input  [7:0]   io_keys_12_2_2,
  input  [7:0]   io_keys_12_2_3,
  input  [7:0]   io_keys_12_3_0,
  input  [7:0]   io_keys_12_3_1,
  input  [7:0]   io_keys_12_3_2,
  input  [7:0]   io_keys_12_3_3,
  input  [7:0]   io_keys_13_0_0,
  input  [7:0]   io_keys_13_0_1,
  input  [7:0]   io_keys_13_0_2,
  input  [7:0]   io_keys_13_0_3,
  input  [7:0]   io_keys_13_1_0,
  input  [7:0]   io_keys_13_1_1,
  input  [7:0]   io_keys_13_1_2,
  input  [7:0]   io_keys_13_1_3,
  input  [7:0]   io_keys_13_2_0,
  input  [7:0]   io_keys_13_2_1,
  input  [7:0]   io_keys_13_2_2,
  input  [7:0]   io_keys_13_2_3,
  input  [7:0]   io_keys_13_3_0,
  input  [7:0]   io_keys_13_3_1,
  input  [7:0]   io_keys_13_3_2,
  input  [7:0]   io_keys_13_3_3,
  input  [7:0]   io_keys_14_0_0,
  input  [7:0]   io_keys_14_0_1,
  input  [7:0]   io_keys_14_0_2,
  input  [7:0]   io_keys_14_0_3,
  input  [7:0]   io_keys_14_1_0,
  input  [7:0]   io_keys_14_1_1,
  input  [7:0]   io_keys_14_1_2,
  input  [7:0]   io_keys_14_1_3,
  input  [7:0]   io_keys_14_2_0,
  input  [7:0]   io_keys_14_2_1,
  input  [7:0]   io_keys_14_2_2,
  input  [7:0]   io_keys_14_2_3,
  input  [7:0]   io_keys_14_3_0,
  input  [7:0]   io_keys_14_3_1,
  input  [7:0]   io_keys_14_3_2,
  input  [7:0]   io_keys_14_3_3,
  input          io_aes256,
  output         io_shiftCyc,
  output         io_shiftRev,
  output         io_shift,
  output         io_ready,
  output [127:0] io_dataOut,
  output [127:0] io_ivOut,
  output         io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] MixColsModule_io_in_0_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_0_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_0_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_0_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_1_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_2_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_in_3_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_0_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_1_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_2_3; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_0; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_1; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_2; // @[AesComponents.scala 91:35]
  wire [7:0] MixColsModule_io_out_3_3; // @[AesComponents.scala 91:35]
  reg [5:0] state; // @[AesDecrypt.scala 53:24]
  wire  _T = state == 6'h0; // @[AesDecrypt.scala 55:25]
  wire  _T_1 = state == 6'h1e; // @[AesDecrypt.scala 55:44]
  reg [127:0] ctSaved; // @[AesDecrypt.scala 62:22]
  reg [7:0] matrix_0_0; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_0_1; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_0_2; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_0_3; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_1_0; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_1_1; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_1_2; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_1_3; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_2_0; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_2_1; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_2_2; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_2_3; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_3_0; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_3_1; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_3_2; // @[AesDecrypt.scala 65:21]
  reg [7:0] matrix_3_3; // @[AesDecrypt.scala 65:21]
  wire [63:0] _T_10 = {matrix_2_0,matrix_2_1,matrix_2_2,matrix_2_3,matrix_3_0,matrix_3_1,matrix_3_2,matrix_3_3}; // @[Cat.scala 29:58]
  wire [63:0] _T_17 = {matrix_0_0,matrix_0_1,matrix_0_2,matrix_0_3,matrix_1_0,matrix_1_1,matrix_1_2,matrix_1_3}; // @[Cat.scala 29:58]
  wire  _T_41 = matrix_0_0[7] ^ matrix_0_0[4]; // @[AesSbox.scala 40:63]
  wire  _T_43 = matrix_0_0[6] ^ matrix_0_0[4]; // @[AesSbox.scala 42:65]
  wire  _T_44 = ~_T_43; // @[AesSbox.scala 42:51]
  wire  _T_46 = matrix_0_0[7] ^ matrix_0_0[6]; // @[AesSbox.scala 42:65]
  wire  _T_47 = ~_T_46; // @[AesSbox.scala 42:51]
  wire  _T_49 = matrix_0_0[4] ^ matrix_0_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_51 = matrix_0_0[3] ^ matrix_0_0[0]; // @[AesSbox.scala 42:65]
  wire  _T_52 = ~_T_51; // @[AesSbox.scala 42:51]
  wire  _T_54 = matrix_0_0[1] ^ matrix_0_0[0]; // @[AesSbox.scala 40:63]
  wire  _T_56 = matrix_0_0[6] ^ _T_41; // @[AesSbox.scala 42:65]
  wire  _T_57 = ~_T_56; // @[AesSbox.scala 42:51]
  wire  _T_59 = _T_44 ^ _T_54; // @[AesSbox.scala 40:63]
  wire  _T_61 = matrix_0_0[0] ^ _T_49; // @[AesSbox.scala 42:65]
  wire  _T_62 = ~_T_61; // @[AesSbox.scala 42:51]
  wire  _T_64 = _T_47 ^ _T_52; // @[AesSbox.scala 40:63]
  wire  _T_66 = _T_47 ^ _T_54; // @[AesSbox.scala 40:63]
  wire  _T_68 = _T_49 ^ _T_54; // @[AesSbox.scala 40:63]
  wire  _T_70 = matrix_0_0[5] ^ _T_49; // @[AesSbox.scala 42:65]
  wire  _T_71 = ~_T_70; // @[AesSbox.scala 42:51]
  wire  _T_73 = matrix_0_0[6] ^ matrix_0_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_75 = matrix_0_0[5] ^ _T_59; // @[AesSbox.scala 42:65]
  wire  _T_76 = ~_T_75; // @[AesSbox.scala 42:51]
  wire  _T_78 = _T_52 ^ _T_73; // @[AesSbox.scala 40:63]
  wire  _T_80 = matrix_0_0[3] ^ _T_57; // @[AesSbox.scala 40:63]
  wire  _T_82 = matrix_0_0[5] ^ matrix_0_0[2]; // @[AesSbox.scala 42:65]
  wire  _T_83 = ~_T_82; // @[AesSbox.scala 42:51]
  wire  _T_85 = matrix_0_0[2] ^ matrix_0_0[1]; // @[AesSbox.scala 42:65]
  wire  _T_86 = ~_T_85; // @[AesSbox.scala 42:51]
  wire  _T_88 = matrix_0_0[5] ^ matrix_0_0[3]; // @[AesSbox.scala 42:65]
  wire  _T_89 = ~_T_88; // @[AesSbox.scala 42:51]
  wire  _T_91 = matrix_0_0[7] ^ _T_83; // @[AesSbox.scala 40:63]
  wire  _T_93 = _T_44 ^ _T_83; // @[AesSbox.scala 40:63]
  wire  _T_95 = _T_73 ^ _T_89; // @[AesSbox.scala 40:63]
  wire  _T_97 = _T_49 ^ _T_86; // @[AesSbox.scala 40:63]
  wire  _T_99 = _T_64 ^ _T_97; // @[AesSbox.scala 40:63]
  wire  _T_101 = _T_64 ^ _T_86; // @[AesSbox.scala 40:63]
  wire  _T_103 = _T_68 ^ _T_95; // @[AesSbox.scala 40:63]
  wire  _T_105 = _T_66 & _T_93; // @[AesSbox.scala 41:63]
  wire  _T_107 = _T_41 & _T_57; // @[AesSbox.scala 41:63]
  wire  _T_109 = _T_101 ^ _T_105; // @[AesSbox.scala 40:63]
  wire  _T_111 = _T_59 & _T_91; // @[AesSbox.scala 41:63]
  wire  _T_113 = _T_111 ^ _T_105; // @[AesSbox.scala 40:63]
  wire  _T_115 = _T_68 & _T_95; // @[AesSbox.scala 41:63]
  wire  _T_117 = _T_44 & _T_62; // @[AesSbox.scala 41:63]
  wire  _T_119 = _T_103 ^ _T_115; // @[AesSbox.scala 40:63]
  wire  _T_121 = _T_78 & _T_76; // @[AesSbox.scala 41:63]
  wire  _T_123 = _T_121 ^ _T_115; // @[AesSbox.scala 40:63]
  wire  _T_125 = _T_49 & _T_99; // @[AesSbox.scala 41:63]
  wire  _T_127 = _T_80 & _T_97; // @[AesSbox.scala 41:63]
  wire  _T_129 = _T_127 ^ _T_125; // @[AesSbox.scala 40:63]
  wire  _T_131 = _T_47 & _T_64; // @[AesSbox.scala 41:63]
  wire  _T_133 = _T_131 ^ _T_125; // @[AesSbox.scala 40:63]
  wire  _T_135 = _T_109 ^ _T_107; // @[AesSbox.scala 40:63]
  wire  _T_137 = _T_113 ^ _T_52; // @[AesSbox.scala 40:63]
  wire  _T_139 = _T_119 ^ _T_117; // @[AesSbox.scala 40:63]
  wire  _T_141 = _T_123 ^ _T_133; // @[AesSbox.scala 40:63]
  wire  _T_143 = _T_135 ^ _T_129; // @[AesSbox.scala 40:63]
  wire  _T_145 = _T_137 ^ _T_133; // @[AesSbox.scala 40:63]
  wire  _T_147 = _T_139 ^ _T_129; // @[AesSbox.scala 40:63]
  wire  _T_149 = _T_141 ^ _T_71; // @[AesSbox.scala 40:63]
  wire  _T_151 = _T_147 ^ _T_149; // @[AesSbox.scala 40:63]
  wire  _T_153 = _T_147 & _T_143; // @[AesSbox.scala 41:63]
  wire  _T_155 = _T_145 ^ _T_153; // @[AesSbox.scala 40:63]
  wire  _T_157 = _T_143 ^ _T_145; // @[AesSbox.scala 40:63]
  wire  _T_159 = _T_149 ^ _T_153; // @[AesSbox.scala 40:63]
  wire  _T_161 = _T_159 & _T_157; // @[AesSbox.scala 41:63]
  wire  _T_163 = _T_155 & _T_151; // @[AesSbox.scala 41:63]
  wire  _T_165 = _T_143 & _T_149; // @[AesSbox.scala 41:63]
  wire  _T_167 = _T_157 & _T_165; // @[AesSbox.scala 41:63]
  wire  _T_169 = _T_157 ^ _T_153; // @[AesSbox.scala 40:63]
  wire  _T_171 = _T_145 & _T_147; // @[AesSbox.scala 41:63]
  wire  _T_173 = _T_151 & _T_171; // @[AesSbox.scala 41:63]
  wire  _T_175 = _T_151 ^ _T_153; // @[AesSbox.scala 40:63]
  wire  _T_177 = _T_145 ^ _T_161; // @[AesSbox.scala 40:63]
  wire  _T_179 = _T_167 ^ _T_169; // @[AesSbox.scala 40:63]
  wire  _T_181 = _T_149 ^ _T_163; // @[AesSbox.scala 40:63]
  wire  _T_183 = _T_173 ^ _T_175; // @[AesSbox.scala 40:63]
  wire  _T_185 = _T_179 ^ _T_183; // @[AesSbox.scala 40:63]
  wire  _T_187 = _T_177 ^ _T_181; // @[AesSbox.scala 40:63]
  wire  _T_189 = _T_177 ^ _T_179; // @[AesSbox.scala 40:63]
  wire  _T_191 = _T_181 ^ _T_183; // @[AesSbox.scala 40:63]
  wire  _T_193 = _T_187 ^ _T_185; // @[AesSbox.scala 40:63]
  wire  _T_195 = _T_191 & _T_93; // @[AesSbox.scala 41:63]
  wire  _T_197 = _T_183 & _T_57; // @[AesSbox.scala 41:63]
  wire  _T_199 = _T_181 & _T_91; // @[AesSbox.scala 41:63]
  wire  _T_201 = _T_189 & _T_95; // @[AesSbox.scala 41:63]
  wire  _T_203 = _T_179 & _T_62; // @[AesSbox.scala 41:63]
  wire  _T_205 = _T_177 & _T_76; // @[AesSbox.scala 41:63]
  wire  _T_207 = _T_187 & _T_99; // @[AesSbox.scala 41:63]
  wire  _T_209 = _T_193 & _T_97; // @[AesSbox.scala 41:63]
  wire  _T_211 = _T_185 & _T_64; // @[AesSbox.scala 41:63]
  wire  _T_213 = _T_191 & _T_66; // @[AesSbox.scala 41:63]
  wire  _T_215 = _T_183 & _T_41; // @[AesSbox.scala 41:63]
  wire  _T_217 = _T_181 & _T_59; // @[AesSbox.scala 41:63]
  wire  _T_219 = _T_189 & _T_68; // @[AesSbox.scala 41:63]
  wire  _T_221 = _T_179 & _T_44; // @[AesSbox.scala 41:63]
  wire  _T_223 = _T_177 & _T_78; // @[AesSbox.scala 41:63]
  wire  _T_225 = _T_187 & _T_49; // @[AesSbox.scala 41:63]
  wire  _T_227 = _T_193 & _T_80; // @[AesSbox.scala 41:63]
  wire  _T_229 = _T_185 & _T_47; // @[AesSbox.scala 41:63]
  wire  _T_231 = _T_207 ^ _T_225; // @[AesSbox.scala 40:63]
  wire  _T_233 = _T_219 ^ _T_221; // @[AesSbox.scala 40:63]
  wire  _T_235 = _T_211 ^ _T_227; // @[AesSbox.scala 40:63]
  wire  _T_237 = _T_197 ^ _T_203; // @[AesSbox.scala 40:63]
  wire  _T_239 = _T_199 ^ _T_215; // @[AesSbox.scala 40:63]
  wire  _T_241 = _T_195 ^ _T_205; // @[AesSbox.scala 40:63]
  wire  _T_243 = _T_201 ^ _T_223; // @[AesSbox.scala 40:63]
  wire  _T_245 = _T_231 ^ _T_233; // @[AesSbox.scala 40:63]
  wire  _T_247 = _T_203 ^ _T_209; // @[AesSbox.scala 40:63]
  wire  _T_249 = _T_213 ^ _T_229; // @[AesSbox.scala 40:63]
  wire  _T_251 = _T_217 ^ _T_239; // @[AesSbox.scala 40:63]
  wire  _T_253 = _T_231 ^ _T_237; // @[AesSbox.scala 40:63]
  wire  _T_255 = _T_195 ^ _T_199; // @[AesSbox.scala 40:63]
  wire  _T_257 = _T_201 ^ _T_205; // @[AesSbox.scala 40:63]
  wire  _T_259 = _T_201 ^ _T_227; // @[AesSbox.scala 40:63]
  wire  _T_261 = _T_211 ^ _T_221; // @[AesSbox.scala 40:63]
  wire  _T_263 = _T_217 ^ _T_225; // @[AesSbox.scala 40:63]
  wire  _T_265 = _T_219 ^ _T_235; // @[AesSbox.scala 40:63]
  wire  _T_267 = _T_229 ^ _T_241; // @[AesSbox.scala 40:63]
  wire  _T_269 = _T_235 ^ _T_237; // @[AesSbox.scala 40:63]
  wire  _T_271 = _T_239 ^ _T_243; // @[AesSbox.scala 40:63]
  wire  _T_273 = _T_235 ^ _T_245; // @[AesSbox.scala 40:63]
  wire  _T_275 = _T_245 ^ _T_247; // @[AesSbox.scala 40:63]
  wire  _T_277 = _T_241 ^ _T_245; // @[AesSbox.scala 40:63]
  wire  _T_279 = _T_243 ^ _T_251; // @[AesSbox.scala 40:63]
  wire  _T_281 = _T_249 ^ _T_253; // @[AesSbox.scala 40:63]
  wire  _T_283 = _T_251 ^ _T_267; // @[AesSbox.scala 40:63]
  wire  _T_285 = _T_253 ^ _T_279; // @[AesSbox.scala 40:63]
  wire  _T_287 = _T_261 ^ _T_271; // @[AesSbox.scala 40:63]
  wire  _T_288 = _T_257 ^ _T_273; // @[AesSbox.scala 40:63]
  wire  _T_289 = _T_281 ^ _T_287; // @[AesSbox.scala 40:63]
  wire  _T_290 = _T_265 ^ _T_285; // @[AesSbox.scala 40:63]
  wire  _T_291 = _T_255 ^ _T_273; // @[AesSbox.scala 40:63]
  wire  _T_292 = _T_275 ^ _T_283; // @[AesSbox.scala 40:63]
  wire  _T_293 = _T_269 ^ _T_277; // @[AesSbox.scala 40:63]
  wire  _T_294 = _T_259 ^ _T_275; // @[AesSbox.scala 40:63]
  wire  _T_295 = _T_249 ^ _T_263; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_0_0 = {_T_288,_T_289,_T_290,_T_291,_T_292,_T_293,_T_294,_T_295}; // @[Cat.scala 29:58]
  wire  _T_320 = matrix_3_1[7] ^ matrix_3_1[4]; // @[AesSbox.scala 40:63]
  wire  _T_322 = matrix_3_1[6] ^ matrix_3_1[4]; // @[AesSbox.scala 42:65]
  wire  _T_323 = ~_T_322; // @[AesSbox.scala 42:51]
  wire  _T_325 = matrix_3_1[7] ^ matrix_3_1[6]; // @[AesSbox.scala 42:65]
  wire  _T_326 = ~_T_325; // @[AesSbox.scala 42:51]
  wire  _T_328 = matrix_3_1[4] ^ matrix_3_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_330 = matrix_3_1[3] ^ matrix_3_1[0]; // @[AesSbox.scala 42:65]
  wire  _T_331 = ~_T_330; // @[AesSbox.scala 42:51]
  wire  _T_333 = matrix_3_1[1] ^ matrix_3_1[0]; // @[AesSbox.scala 40:63]
  wire  _T_335 = matrix_3_1[6] ^ _T_320; // @[AesSbox.scala 42:65]
  wire  _T_336 = ~_T_335; // @[AesSbox.scala 42:51]
  wire  _T_338 = _T_323 ^ _T_333; // @[AesSbox.scala 40:63]
  wire  _T_340 = matrix_3_1[0] ^ _T_328; // @[AesSbox.scala 42:65]
  wire  _T_341 = ~_T_340; // @[AesSbox.scala 42:51]
  wire  _T_343 = _T_326 ^ _T_331; // @[AesSbox.scala 40:63]
  wire  _T_345 = _T_326 ^ _T_333; // @[AesSbox.scala 40:63]
  wire  _T_347 = _T_328 ^ _T_333; // @[AesSbox.scala 40:63]
  wire  _T_349 = matrix_3_1[5] ^ _T_328; // @[AesSbox.scala 42:65]
  wire  _T_350 = ~_T_349; // @[AesSbox.scala 42:51]
  wire  _T_352 = matrix_3_1[6] ^ matrix_3_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_354 = matrix_3_1[5] ^ _T_338; // @[AesSbox.scala 42:65]
  wire  _T_355 = ~_T_354; // @[AesSbox.scala 42:51]
  wire  _T_357 = _T_331 ^ _T_352; // @[AesSbox.scala 40:63]
  wire  _T_359 = matrix_3_1[3] ^ _T_336; // @[AesSbox.scala 40:63]
  wire  _T_361 = matrix_3_1[5] ^ matrix_3_1[2]; // @[AesSbox.scala 42:65]
  wire  _T_362 = ~_T_361; // @[AesSbox.scala 42:51]
  wire  _T_364 = matrix_3_1[2] ^ matrix_3_1[1]; // @[AesSbox.scala 42:65]
  wire  _T_365 = ~_T_364; // @[AesSbox.scala 42:51]
  wire  _T_367 = matrix_3_1[5] ^ matrix_3_1[3]; // @[AesSbox.scala 42:65]
  wire  _T_368 = ~_T_367; // @[AesSbox.scala 42:51]
  wire  _T_370 = matrix_3_1[7] ^ _T_362; // @[AesSbox.scala 40:63]
  wire  _T_372 = _T_323 ^ _T_362; // @[AesSbox.scala 40:63]
  wire  _T_374 = _T_352 ^ _T_368; // @[AesSbox.scala 40:63]
  wire  _T_376 = _T_328 ^ _T_365; // @[AesSbox.scala 40:63]
  wire  _T_378 = _T_343 ^ _T_376; // @[AesSbox.scala 40:63]
  wire  _T_380 = _T_343 ^ _T_365; // @[AesSbox.scala 40:63]
  wire  _T_382 = _T_347 ^ _T_374; // @[AesSbox.scala 40:63]
  wire  _T_384 = _T_345 & _T_372; // @[AesSbox.scala 41:63]
  wire  _T_386 = _T_320 & _T_336; // @[AesSbox.scala 41:63]
  wire  _T_388 = _T_380 ^ _T_384; // @[AesSbox.scala 40:63]
  wire  _T_390 = _T_338 & _T_370; // @[AesSbox.scala 41:63]
  wire  _T_392 = _T_390 ^ _T_384; // @[AesSbox.scala 40:63]
  wire  _T_394 = _T_347 & _T_374; // @[AesSbox.scala 41:63]
  wire  _T_396 = _T_323 & _T_341; // @[AesSbox.scala 41:63]
  wire  _T_398 = _T_382 ^ _T_394; // @[AesSbox.scala 40:63]
  wire  _T_400 = _T_357 & _T_355; // @[AesSbox.scala 41:63]
  wire  _T_402 = _T_400 ^ _T_394; // @[AesSbox.scala 40:63]
  wire  _T_404 = _T_328 & _T_378; // @[AesSbox.scala 41:63]
  wire  _T_406 = _T_359 & _T_376; // @[AesSbox.scala 41:63]
  wire  _T_408 = _T_406 ^ _T_404; // @[AesSbox.scala 40:63]
  wire  _T_410 = _T_326 & _T_343; // @[AesSbox.scala 41:63]
  wire  _T_412 = _T_410 ^ _T_404; // @[AesSbox.scala 40:63]
  wire  _T_414 = _T_388 ^ _T_386; // @[AesSbox.scala 40:63]
  wire  _T_416 = _T_392 ^ _T_331; // @[AesSbox.scala 40:63]
  wire  _T_418 = _T_398 ^ _T_396; // @[AesSbox.scala 40:63]
  wire  _T_420 = _T_402 ^ _T_412; // @[AesSbox.scala 40:63]
  wire  _T_422 = _T_414 ^ _T_408; // @[AesSbox.scala 40:63]
  wire  _T_424 = _T_416 ^ _T_412; // @[AesSbox.scala 40:63]
  wire  _T_426 = _T_418 ^ _T_408; // @[AesSbox.scala 40:63]
  wire  _T_428 = _T_420 ^ _T_350; // @[AesSbox.scala 40:63]
  wire  _T_430 = _T_426 ^ _T_428; // @[AesSbox.scala 40:63]
  wire  _T_432 = _T_426 & _T_422; // @[AesSbox.scala 41:63]
  wire  _T_434 = _T_424 ^ _T_432; // @[AesSbox.scala 40:63]
  wire  _T_436 = _T_422 ^ _T_424; // @[AesSbox.scala 40:63]
  wire  _T_438 = _T_428 ^ _T_432; // @[AesSbox.scala 40:63]
  wire  _T_440 = _T_438 & _T_436; // @[AesSbox.scala 41:63]
  wire  _T_442 = _T_434 & _T_430; // @[AesSbox.scala 41:63]
  wire  _T_444 = _T_422 & _T_428; // @[AesSbox.scala 41:63]
  wire  _T_446 = _T_436 & _T_444; // @[AesSbox.scala 41:63]
  wire  _T_448 = _T_436 ^ _T_432; // @[AesSbox.scala 40:63]
  wire  _T_450 = _T_424 & _T_426; // @[AesSbox.scala 41:63]
  wire  _T_452 = _T_430 & _T_450; // @[AesSbox.scala 41:63]
  wire  _T_454 = _T_430 ^ _T_432; // @[AesSbox.scala 40:63]
  wire  _T_456 = _T_424 ^ _T_440; // @[AesSbox.scala 40:63]
  wire  _T_458 = _T_446 ^ _T_448; // @[AesSbox.scala 40:63]
  wire  _T_460 = _T_428 ^ _T_442; // @[AesSbox.scala 40:63]
  wire  _T_462 = _T_452 ^ _T_454; // @[AesSbox.scala 40:63]
  wire  _T_464 = _T_458 ^ _T_462; // @[AesSbox.scala 40:63]
  wire  _T_466 = _T_456 ^ _T_460; // @[AesSbox.scala 40:63]
  wire  _T_468 = _T_456 ^ _T_458; // @[AesSbox.scala 40:63]
  wire  _T_470 = _T_460 ^ _T_462; // @[AesSbox.scala 40:63]
  wire  _T_472 = _T_466 ^ _T_464; // @[AesSbox.scala 40:63]
  wire  _T_474 = _T_470 & _T_372; // @[AesSbox.scala 41:63]
  wire  _T_476 = _T_462 & _T_336; // @[AesSbox.scala 41:63]
  wire  _T_478 = _T_460 & _T_370; // @[AesSbox.scala 41:63]
  wire  _T_480 = _T_468 & _T_374; // @[AesSbox.scala 41:63]
  wire  _T_482 = _T_458 & _T_341; // @[AesSbox.scala 41:63]
  wire  _T_484 = _T_456 & _T_355; // @[AesSbox.scala 41:63]
  wire  _T_486 = _T_466 & _T_378; // @[AesSbox.scala 41:63]
  wire  _T_488 = _T_472 & _T_376; // @[AesSbox.scala 41:63]
  wire  _T_490 = _T_464 & _T_343; // @[AesSbox.scala 41:63]
  wire  _T_492 = _T_470 & _T_345; // @[AesSbox.scala 41:63]
  wire  _T_494 = _T_462 & _T_320; // @[AesSbox.scala 41:63]
  wire  _T_496 = _T_460 & _T_338; // @[AesSbox.scala 41:63]
  wire  _T_498 = _T_468 & _T_347; // @[AesSbox.scala 41:63]
  wire  _T_500 = _T_458 & _T_323; // @[AesSbox.scala 41:63]
  wire  _T_502 = _T_456 & _T_357; // @[AesSbox.scala 41:63]
  wire  _T_504 = _T_466 & _T_328; // @[AesSbox.scala 41:63]
  wire  _T_506 = _T_472 & _T_359; // @[AesSbox.scala 41:63]
  wire  _T_508 = _T_464 & _T_326; // @[AesSbox.scala 41:63]
  wire  _T_510 = _T_486 ^ _T_504; // @[AesSbox.scala 40:63]
  wire  _T_512 = _T_498 ^ _T_500; // @[AesSbox.scala 40:63]
  wire  _T_514 = _T_490 ^ _T_506; // @[AesSbox.scala 40:63]
  wire  _T_516 = _T_476 ^ _T_482; // @[AesSbox.scala 40:63]
  wire  _T_518 = _T_478 ^ _T_494; // @[AesSbox.scala 40:63]
  wire  _T_520 = _T_474 ^ _T_484; // @[AesSbox.scala 40:63]
  wire  _T_522 = _T_480 ^ _T_502; // @[AesSbox.scala 40:63]
  wire  _T_524 = _T_510 ^ _T_512; // @[AesSbox.scala 40:63]
  wire  _T_526 = _T_482 ^ _T_488; // @[AesSbox.scala 40:63]
  wire  _T_528 = _T_492 ^ _T_508; // @[AesSbox.scala 40:63]
  wire  _T_530 = _T_496 ^ _T_518; // @[AesSbox.scala 40:63]
  wire  _T_532 = _T_510 ^ _T_516; // @[AesSbox.scala 40:63]
  wire  _T_534 = _T_474 ^ _T_478; // @[AesSbox.scala 40:63]
  wire  _T_536 = _T_480 ^ _T_484; // @[AesSbox.scala 40:63]
  wire  _T_538 = _T_480 ^ _T_506; // @[AesSbox.scala 40:63]
  wire  _T_540 = _T_490 ^ _T_500; // @[AesSbox.scala 40:63]
  wire  _T_542 = _T_496 ^ _T_504; // @[AesSbox.scala 40:63]
  wire  _T_544 = _T_498 ^ _T_514; // @[AesSbox.scala 40:63]
  wire  _T_546 = _T_508 ^ _T_520; // @[AesSbox.scala 40:63]
  wire  _T_548 = _T_514 ^ _T_516; // @[AesSbox.scala 40:63]
  wire  _T_550 = _T_518 ^ _T_522; // @[AesSbox.scala 40:63]
  wire  _T_552 = _T_514 ^ _T_524; // @[AesSbox.scala 40:63]
  wire  _T_554 = _T_524 ^ _T_526; // @[AesSbox.scala 40:63]
  wire  _T_556 = _T_520 ^ _T_524; // @[AesSbox.scala 40:63]
  wire  _T_558 = _T_522 ^ _T_530; // @[AesSbox.scala 40:63]
  wire  _T_560 = _T_528 ^ _T_532; // @[AesSbox.scala 40:63]
  wire  _T_562 = _T_530 ^ _T_546; // @[AesSbox.scala 40:63]
  wire  _T_564 = _T_532 ^ _T_558; // @[AesSbox.scala 40:63]
  wire  _T_566 = _T_540 ^ _T_550; // @[AesSbox.scala 40:63]
  wire  _T_567 = _T_536 ^ _T_552; // @[AesSbox.scala 40:63]
  wire  _T_568 = _T_560 ^ _T_566; // @[AesSbox.scala 40:63]
  wire  _T_569 = _T_544 ^ _T_564; // @[AesSbox.scala 40:63]
  wire  _T_570 = _T_534 ^ _T_552; // @[AesSbox.scala 40:63]
  wire  _T_571 = _T_554 ^ _T_562; // @[AesSbox.scala 40:63]
  wire  _T_572 = _T_548 ^ _T_556; // @[AesSbox.scala 40:63]
  wire  _T_573 = _T_538 ^ _T_554; // @[AesSbox.scala 40:63]
  wire  _T_574 = _T_528 ^ _T_542; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_0_1 = {_T_567,_T_568,_T_569,_T_570,_T_571,_T_572,_T_573,_T_574}; // @[Cat.scala 29:58]
  wire  _T_599 = matrix_2_2[7] ^ matrix_2_2[4]; // @[AesSbox.scala 40:63]
  wire  _T_601 = matrix_2_2[6] ^ matrix_2_2[4]; // @[AesSbox.scala 42:65]
  wire  _T_602 = ~_T_601; // @[AesSbox.scala 42:51]
  wire  _T_604 = matrix_2_2[7] ^ matrix_2_2[6]; // @[AesSbox.scala 42:65]
  wire  _T_605 = ~_T_604; // @[AesSbox.scala 42:51]
  wire  _T_607 = matrix_2_2[4] ^ matrix_2_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_609 = matrix_2_2[3] ^ matrix_2_2[0]; // @[AesSbox.scala 42:65]
  wire  _T_610 = ~_T_609; // @[AesSbox.scala 42:51]
  wire  _T_612 = matrix_2_2[1] ^ matrix_2_2[0]; // @[AesSbox.scala 40:63]
  wire  _T_614 = matrix_2_2[6] ^ _T_599; // @[AesSbox.scala 42:65]
  wire  _T_615 = ~_T_614; // @[AesSbox.scala 42:51]
  wire  _T_617 = _T_602 ^ _T_612; // @[AesSbox.scala 40:63]
  wire  _T_619 = matrix_2_2[0] ^ _T_607; // @[AesSbox.scala 42:65]
  wire  _T_620 = ~_T_619; // @[AesSbox.scala 42:51]
  wire  _T_622 = _T_605 ^ _T_610; // @[AesSbox.scala 40:63]
  wire  _T_624 = _T_605 ^ _T_612; // @[AesSbox.scala 40:63]
  wire  _T_626 = _T_607 ^ _T_612; // @[AesSbox.scala 40:63]
  wire  _T_628 = matrix_2_2[5] ^ _T_607; // @[AesSbox.scala 42:65]
  wire  _T_629 = ~_T_628; // @[AesSbox.scala 42:51]
  wire  _T_631 = matrix_2_2[6] ^ matrix_2_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_633 = matrix_2_2[5] ^ _T_617; // @[AesSbox.scala 42:65]
  wire  _T_634 = ~_T_633; // @[AesSbox.scala 42:51]
  wire  _T_636 = _T_610 ^ _T_631; // @[AesSbox.scala 40:63]
  wire  _T_638 = matrix_2_2[3] ^ _T_615; // @[AesSbox.scala 40:63]
  wire  _T_640 = matrix_2_2[5] ^ matrix_2_2[2]; // @[AesSbox.scala 42:65]
  wire  _T_641 = ~_T_640; // @[AesSbox.scala 42:51]
  wire  _T_643 = matrix_2_2[2] ^ matrix_2_2[1]; // @[AesSbox.scala 42:65]
  wire  _T_644 = ~_T_643; // @[AesSbox.scala 42:51]
  wire  _T_646 = matrix_2_2[5] ^ matrix_2_2[3]; // @[AesSbox.scala 42:65]
  wire  _T_647 = ~_T_646; // @[AesSbox.scala 42:51]
  wire  _T_649 = matrix_2_2[7] ^ _T_641; // @[AesSbox.scala 40:63]
  wire  _T_651 = _T_602 ^ _T_641; // @[AesSbox.scala 40:63]
  wire  _T_653 = _T_631 ^ _T_647; // @[AesSbox.scala 40:63]
  wire  _T_655 = _T_607 ^ _T_644; // @[AesSbox.scala 40:63]
  wire  _T_657 = _T_622 ^ _T_655; // @[AesSbox.scala 40:63]
  wire  _T_659 = _T_622 ^ _T_644; // @[AesSbox.scala 40:63]
  wire  _T_661 = _T_626 ^ _T_653; // @[AesSbox.scala 40:63]
  wire  _T_663 = _T_624 & _T_651; // @[AesSbox.scala 41:63]
  wire  _T_665 = _T_599 & _T_615; // @[AesSbox.scala 41:63]
  wire  _T_667 = _T_659 ^ _T_663; // @[AesSbox.scala 40:63]
  wire  _T_669 = _T_617 & _T_649; // @[AesSbox.scala 41:63]
  wire  _T_671 = _T_669 ^ _T_663; // @[AesSbox.scala 40:63]
  wire  _T_673 = _T_626 & _T_653; // @[AesSbox.scala 41:63]
  wire  _T_675 = _T_602 & _T_620; // @[AesSbox.scala 41:63]
  wire  _T_677 = _T_661 ^ _T_673; // @[AesSbox.scala 40:63]
  wire  _T_679 = _T_636 & _T_634; // @[AesSbox.scala 41:63]
  wire  _T_681 = _T_679 ^ _T_673; // @[AesSbox.scala 40:63]
  wire  _T_683 = _T_607 & _T_657; // @[AesSbox.scala 41:63]
  wire  _T_685 = _T_638 & _T_655; // @[AesSbox.scala 41:63]
  wire  _T_687 = _T_685 ^ _T_683; // @[AesSbox.scala 40:63]
  wire  _T_689 = _T_605 & _T_622; // @[AesSbox.scala 41:63]
  wire  _T_691 = _T_689 ^ _T_683; // @[AesSbox.scala 40:63]
  wire  _T_693 = _T_667 ^ _T_665; // @[AesSbox.scala 40:63]
  wire  _T_695 = _T_671 ^ _T_610; // @[AesSbox.scala 40:63]
  wire  _T_697 = _T_677 ^ _T_675; // @[AesSbox.scala 40:63]
  wire  _T_699 = _T_681 ^ _T_691; // @[AesSbox.scala 40:63]
  wire  _T_701 = _T_693 ^ _T_687; // @[AesSbox.scala 40:63]
  wire  _T_703 = _T_695 ^ _T_691; // @[AesSbox.scala 40:63]
  wire  _T_705 = _T_697 ^ _T_687; // @[AesSbox.scala 40:63]
  wire  _T_707 = _T_699 ^ _T_629; // @[AesSbox.scala 40:63]
  wire  _T_709 = _T_705 ^ _T_707; // @[AesSbox.scala 40:63]
  wire  _T_711 = _T_705 & _T_701; // @[AesSbox.scala 41:63]
  wire  _T_713 = _T_703 ^ _T_711; // @[AesSbox.scala 40:63]
  wire  _T_715 = _T_701 ^ _T_703; // @[AesSbox.scala 40:63]
  wire  _T_717 = _T_707 ^ _T_711; // @[AesSbox.scala 40:63]
  wire  _T_719 = _T_717 & _T_715; // @[AesSbox.scala 41:63]
  wire  _T_721 = _T_713 & _T_709; // @[AesSbox.scala 41:63]
  wire  _T_723 = _T_701 & _T_707; // @[AesSbox.scala 41:63]
  wire  _T_725 = _T_715 & _T_723; // @[AesSbox.scala 41:63]
  wire  _T_727 = _T_715 ^ _T_711; // @[AesSbox.scala 40:63]
  wire  _T_729 = _T_703 & _T_705; // @[AesSbox.scala 41:63]
  wire  _T_731 = _T_709 & _T_729; // @[AesSbox.scala 41:63]
  wire  _T_733 = _T_709 ^ _T_711; // @[AesSbox.scala 40:63]
  wire  _T_735 = _T_703 ^ _T_719; // @[AesSbox.scala 40:63]
  wire  _T_737 = _T_725 ^ _T_727; // @[AesSbox.scala 40:63]
  wire  _T_739 = _T_707 ^ _T_721; // @[AesSbox.scala 40:63]
  wire  _T_741 = _T_731 ^ _T_733; // @[AesSbox.scala 40:63]
  wire  _T_743 = _T_737 ^ _T_741; // @[AesSbox.scala 40:63]
  wire  _T_745 = _T_735 ^ _T_739; // @[AesSbox.scala 40:63]
  wire  _T_747 = _T_735 ^ _T_737; // @[AesSbox.scala 40:63]
  wire  _T_749 = _T_739 ^ _T_741; // @[AesSbox.scala 40:63]
  wire  _T_751 = _T_745 ^ _T_743; // @[AesSbox.scala 40:63]
  wire  _T_753 = _T_749 & _T_651; // @[AesSbox.scala 41:63]
  wire  _T_755 = _T_741 & _T_615; // @[AesSbox.scala 41:63]
  wire  _T_757 = _T_739 & _T_649; // @[AesSbox.scala 41:63]
  wire  _T_759 = _T_747 & _T_653; // @[AesSbox.scala 41:63]
  wire  _T_761 = _T_737 & _T_620; // @[AesSbox.scala 41:63]
  wire  _T_763 = _T_735 & _T_634; // @[AesSbox.scala 41:63]
  wire  _T_765 = _T_745 & _T_657; // @[AesSbox.scala 41:63]
  wire  _T_767 = _T_751 & _T_655; // @[AesSbox.scala 41:63]
  wire  _T_769 = _T_743 & _T_622; // @[AesSbox.scala 41:63]
  wire  _T_771 = _T_749 & _T_624; // @[AesSbox.scala 41:63]
  wire  _T_773 = _T_741 & _T_599; // @[AesSbox.scala 41:63]
  wire  _T_775 = _T_739 & _T_617; // @[AesSbox.scala 41:63]
  wire  _T_777 = _T_747 & _T_626; // @[AesSbox.scala 41:63]
  wire  _T_779 = _T_737 & _T_602; // @[AesSbox.scala 41:63]
  wire  _T_781 = _T_735 & _T_636; // @[AesSbox.scala 41:63]
  wire  _T_783 = _T_745 & _T_607; // @[AesSbox.scala 41:63]
  wire  _T_785 = _T_751 & _T_638; // @[AesSbox.scala 41:63]
  wire  _T_787 = _T_743 & _T_605; // @[AesSbox.scala 41:63]
  wire  _T_789 = _T_765 ^ _T_783; // @[AesSbox.scala 40:63]
  wire  _T_791 = _T_777 ^ _T_779; // @[AesSbox.scala 40:63]
  wire  _T_793 = _T_769 ^ _T_785; // @[AesSbox.scala 40:63]
  wire  _T_795 = _T_755 ^ _T_761; // @[AesSbox.scala 40:63]
  wire  _T_797 = _T_757 ^ _T_773; // @[AesSbox.scala 40:63]
  wire  _T_799 = _T_753 ^ _T_763; // @[AesSbox.scala 40:63]
  wire  _T_801 = _T_759 ^ _T_781; // @[AesSbox.scala 40:63]
  wire  _T_803 = _T_789 ^ _T_791; // @[AesSbox.scala 40:63]
  wire  _T_805 = _T_761 ^ _T_767; // @[AesSbox.scala 40:63]
  wire  _T_807 = _T_771 ^ _T_787; // @[AesSbox.scala 40:63]
  wire  _T_809 = _T_775 ^ _T_797; // @[AesSbox.scala 40:63]
  wire  _T_811 = _T_789 ^ _T_795; // @[AesSbox.scala 40:63]
  wire  _T_813 = _T_753 ^ _T_757; // @[AesSbox.scala 40:63]
  wire  _T_815 = _T_759 ^ _T_763; // @[AesSbox.scala 40:63]
  wire  _T_817 = _T_759 ^ _T_785; // @[AesSbox.scala 40:63]
  wire  _T_819 = _T_769 ^ _T_779; // @[AesSbox.scala 40:63]
  wire  _T_821 = _T_775 ^ _T_783; // @[AesSbox.scala 40:63]
  wire  _T_823 = _T_777 ^ _T_793; // @[AesSbox.scala 40:63]
  wire  _T_825 = _T_787 ^ _T_799; // @[AesSbox.scala 40:63]
  wire  _T_827 = _T_793 ^ _T_795; // @[AesSbox.scala 40:63]
  wire  _T_829 = _T_797 ^ _T_801; // @[AesSbox.scala 40:63]
  wire  _T_831 = _T_793 ^ _T_803; // @[AesSbox.scala 40:63]
  wire  _T_833 = _T_803 ^ _T_805; // @[AesSbox.scala 40:63]
  wire  _T_835 = _T_799 ^ _T_803; // @[AesSbox.scala 40:63]
  wire  _T_837 = _T_801 ^ _T_809; // @[AesSbox.scala 40:63]
  wire  _T_839 = _T_807 ^ _T_811; // @[AesSbox.scala 40:63]
  wire  _T_841 = _T_809 ^ _T_825; // @[AesSbox.scala 40:63]
  wire  _T_843 = _T_811 ^ _T_837; // @[AesSbox.scala 40:63]
  wire  _T_845 = _T_819 ^ _T_829; // @[AesSbox.scala 40:63]
  wire  _T_846 = _T_815 ^ _T_831; // @[AesSbox.scala 40:63]
  wire  _T_847 = _T_839 ^ _T_845; // @[AesSbox.scala 40:63]
  wire  _T_848 = _T_823 ^ _T_843; // @[AesSbox.scala 40:63]
  wire  _T_849 = _T_813 ^ _T_831; // @[AesSbox.scala 40:63]
  wire  _T_850 = _T_833 ^ _T_841; // @[AesSbox.scala 40:63]
  wire  _T_851 = _T_827 ^ _T_835; // @[AesSbox.scala 40:63]
  wire  _T_852 = _T_817 ^ _T_833; // @[AesSbox.scala 40:63]
  wire  _T_853 = _T_807 ^ _T_821; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_0_2 = {_T_846,_T_847,_T_848,_T_849,_T_850,_T_851,_T_852,_T_853}; // @[Cat.scala 29:58]
  wire  _T_878 = matrix_1_3[7] ^ matrix_1_3[4]; // @[AesSbox.scala 40:63]
  wire  _T_880 = matrix_1_3[6] ^ matrix_1_3[4]; // @[AesSbox.scala 42:65]
  wire  _T_881 = ~_T_880; // @[AesSbox.scala 42:51]
  wire  _T_883 = matrix_1_3[7] ^ matrix_1_3[6]; // @[AesSbox.scala 42:65]
  wire  _T_884 = ~_T_883; // @[AesSbox.scala 42:51]
  wire  _T_886 = matrix_1_3[4] ^ matrix_1_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_888 = matrix_1_3[3] ^ matrix_1_3[0]; // @[AesSbox.scala 42:65]
  wire  _T_889 = ~_T_888; // @[AesSbox.scala 42:51]
  wire  _T_891 = matrix_1_3[1] ^ matrix_1_3[0]; // @[AesSbox.scala 40:63]
  wire  _T_893 = matrix_1_3[6] ^ _T_878; // @[AesSbox.scala 42:65]
  wire  _T_894 = ~_T_893; // @[AesSbox.scala 42:51]
  wire  _T_896 = _T_881 ^ _T_891; // @[AesSbox.scala 40:63]
  wire  _T_898 = matrix_1_3[0] ^ _T_886; // @[AesSbox.scala 42:65]
  wire  _T_899 = ~_T_898; // @[AesSbox.scala 42:51]
  wire  _T_901 = _T_884 ^ _T_889; // @[AesSbox.scala 40:63]
  wire  _T_903 = _T_884 ^ _T_891; // @[AesSbox.scala 40:63]
  wire  _T_905 = _T_886 ^ _T_891; // @[AesSbox.scala 40:63]
  wire  _T_907 = matrix_1_3[5] ^ _T_886; // @[AesSbox.scala 42:65]
  wire  _T_908 = ~_T_907; // @[AesSbox.scala 42:51]
  wire  _T_910 = matrix_1_3[6] ^ matrix_1_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_912 = matrix_1_3[5] ^ _T_896; // @[AesSbox.scala 42:65]
  wire  _T_913 = ~_T_912; // @[AesSbox.scala 42:51]
  wire  _T_915 = _T_889 ^ _T_910; // @[AesSbox.scala 40:63]
  wire  _T_917 = matrix_1_3[3] ^ _T_894; // @[AesSbox.scala 40:63]
  wire  _T_919 = matrix_1_3[5] ^ matrix_1_3[2]; // @[AesSbox.scala 42:65]
  wire  _T_920 = ~_T_919; // @[AesSbox.scala 42:51]
  wire  _T_922 = matrix_1_3[2] ^ matrix_1_3[1]; // @[AesSbox.scala 42:65]
  wire  _T_923 = ~_T_922; // @[AesSbox.scala 42:51]
  wire  _T_925 = matrix_1_3[5] ^ matrix_1_3[3]; // @[AesSbox.scala 42:65]
  wire  _T_926 = ~_T_925; // @[AesSbox.scala 42:51]
  wire  _T_928 = matrix_1_3[7] ^ _T_920; // @[AesSbox.scala 40:63]
  wire  _T_930 = _T_881 ^ _T_920; // @[AesSbox.scala 40:63]
  wire  _T_932 = _T_910 ^ _T_926; // @[AesSbox.scala 40:63]
  wire  _T_934 = _T_886 ^ _T_923; // @[AesSbox.scala 40:63]
  wire  _T_936 = _T_901 ^ _T_934; // @[AesSbox.scala 40:63]
  wire  _T_938 = _T_901 ^ _T_923; // @[AesSbox.scala 40:63]
  wire  _T_940 = _T_905 ^ _T_932; // @[AesSbox.scala 40:63]
  wire  _T_942 = _T_903 & _T_930; // @[AesSbox.scala 41:63]
  wire  _T_944 = _T_878 & _T_894; // @[AesSbox.scala 41:63]
  wire  _T_946 = _T_938 ^ _T_942; // @[AesSbox.scala 40:63]
  wire  _T_948 = _T_896 & _T_928; // @[AesSbox.scala 41:63]
  wire  _T_950 = _T_948 ^ _T_942; // @[AesSbox.scala 40:63]
  wire  _T_952 = _T_905 & _T_932; // @[AesSbox.scala 41:63]
  wire  _T_954 = _T_881 & _T_899; // @[AesSbox.scala 41:63]
  wire  _T_956 = _T_940 ^ _T_952; // @[AesSbox.scala 40:63]
  wire  _T_958 = _T_915 & _T_913; // @[AesSbox.scala 41:63]
  wire  _T_960 = _T_958 ^ _T_952; // @[AesSbox.scala 40:63]
  wire  _T_962 = _T_886 & _T_936; // @[AesSbox.scala 41:63]
  wire  _T_964 = _T_917 & _T_934; // @[AesSbox.scala 41:63]
  wire  _T_966 = _T_964 ^ _T_962; // @[AesSbox.scala 40:63]
  wire  _T_968 = _T_884 & _T_901; // @[AesSbox.scala 41:63]
  wire  _T_970 = _T_968 ^ _T_962; // @[AesSbox.scala 40:63]
  wire  _T_972 = _T_946 ^ _T_944; // @[AesSbox.scala 40:63]
  wire  _T_974 = _T_950 ^ _T_889; // @[AesSbox.scala 40:63]
  wire  _T_976 = _T_956 ^ _T_954; // @[AesSbox.scala 40:63]
  wire  _T_978 = _T_960 ^ _T_970; // @[AesSbox.scala 40:63]
  wire  _T_980 = _T_972 ^ _T_966; // @[AesSbox.scala 40:63]
  wire  _T_982 = _T_974 ^ _T_970; // @[AesSbox.scala 40:63]
  wire  _T_984 = _T_976 ^ _T_966; // @[AesSbox.scala 40:63]
  wire  _T_986 = _T_978 ^ _T_908; // @[AesSbox.scala 40:63]
  wire  _T_988 = _T_984 ^ _T_986; // @[AesSbox.scala 40:63]
  wire  _T_990 = _T_984 & _T_980; // @[AesSbox.scala 41:63]
  wire  _T_992 = _T_982 ^ _T_990; // @[AesSbox.scala 40:63]
  wire  _T_994 = _T_980 ^ _T_982; // @[AesSbox.scala 40:63]
  wire  _T_996 = _T_986 ^ _T_990; // @[AesSbox.scala 40:63]
  wire  _T_998 = _T_996 & _T_994; // @[AesSbox.scala 41:63]
  wire  _T_1000 = _T_992 & _T_988; // @[AesSbox.scala 41:63]
  wire  _T_1002 = _T_980 & _T_986; // @[AesSbox.scala 41:63]
  wire  _T_1004 = _T_994 & _T_1002; // @[AesSbox.scala 41:63]
  wire  _T_1006 = _T_994 ^ _T_990; // @[AesSbox.scala 40:63]
  wire  _T_1008 = _T_982 & _T_984; // @[AesSbox.scala 41:63]
  wire  _T_1010 = _T_988 & _T_1008; // @[AesSbox.scala 41:63]
  wire  _T_1012 = _T_988 ^ _T_990; // @[AesSbox.scala 40:63]
  wire  _T_1014 = _T_982 ^ _T_998; // @[AesSbox.scala 40:63]
  wire  _T_1016 = _T_1004 ^ _T_1006; // @[AesSbox.scala 40:63]
  wire  _T_1018 = _T_986 ^ _T_1000; // @[AesSbox.scala 40:63]
  wire  _T_1020 = _T_1010 ^ _T_1012; // @[AesSbox.scala 40:63]
  wire  _T_1022 = _T_1016 ^ _T_1020; // @[AesSbox.scala 40:63]
  wire  _T_1024 = _T_1014 ^ _T_1018; // @[AesSbox.scala 40:63]
  wire  _T_1026 = _T_1014 ^ _T_1016; // @[AesSbox.scala 40:63]
  wire  _T_1028 = _T_1018 ^ _T_1020; // @[AesSbox.scala 40:63]
  wire  _T_1030 = _T_1024 ^ _T_1022; // @[AesSbox.scala 40:63]
  wire  _T_1032 = _T_1028 & _T_930; // @[AesSbox.scala 41:63]
  wire  _T_1034 = _T_1020 & _T_894; // @[AesSbox.scala 41:63]
  wire  _T_1036 = _T_1018 & _T_928; // @[AesSbox.scala 41:63]
  wire  _T_1038 = _T_1026 & _T_932; // @[AesSbox.scala 41:63]
  wire  _T_1040 = _T_1016 & _T_899; // @[AesSbox.scala 41:63]
  wire  _T_1042 = _T_1014 & _T_913; // @[AesSbox.scala 41:63]
  wire  _T_1044 = _T_1024 & _T_936; // @[AesSbox.scala 41:63]
  wire  _T_1046 = _T_1030 & _T_934; // @[AesSbox.scala 41:63]
  wire  _T_1048 = _T_1022 & _T_901; // @[AesSbox.scala 41:63]
  wire  _T_1050 = _T_1028 & _T_903; // @[AesSbox.scala 41:63]
  wire  _T_1052 = _T_1020 & _T_878; // @[AesSbox.scala 41:63]
  wire  _T_1054 = _T_1018 & _T_896; // @[AesSbox.scala 41:63]
  wire  _T_1056 = _T_1026 & _T_905; // @[AesSbox.scala 41:63]
  wire  _T_1058 = _T_1016 & _T_881; // @[AesSbox.scala 41:63]
  wire  _T_1060 = _T_1014 & _T_915; // @[AesSbox.scala 41:63]
  wire  _T_1062 = _T_1024 & _T_886; // @[AesSbox.scala 41:63]
  wire  _T_1064 = _T_1030 & _T_917; // @[AesSbox.scala 41:63]
  wire  _T_1066 = _T_1022 & _T_884; // @[AesSbox.scala 41:63]
  wire  _T_1068 = _T_1044 ^ _T_1062; // @[AesSbox.scala 40:63]
  wire  _T_1070 = _T_1056 ^ _T_1058; // @[AesSbox.scala 40:63]
  wire  _T_1072 = _T_1048 ^ _T_1064; // @[AesSbox.scala 40:63]
  wire  _T_1074 = _T_1034 ^ _T_1040; // @[AesSbox.scala 40:63]
  wire  _T_1076 = _T_1036 ^ _T_1052; // @[AesSbox.scala 40:63]
  wire  _T_1078 = _T_1032 ^ _T_1042; // @[AesSbox.scala 40:63]
  wire  _T_1080 = _T_1038 ^ _T_1060; // @[AesSbox.scala 40:63]
  wire  _T_1082 = _T_1068 ^ _T_1070; // @[AesSbox.scala 40:63]
  wire  _T_1084 = _T_1040 ^ _T_1046; // @[AesSbox.scala 40:63]
  wire  _T_1086 = _T_1050 ^ _T_1066; // @[AesSbox.scala 40:63]
  wire  _T_1088 = _T_1054 ^ _T_1076; // @[AesSbox.scala 40:63]
  wire  _T_1090 = _T_1068 ^ _T_1074; // @[AesSbox.scala 40:63]
  wire  _T_1092 = _T_1032 ^ _T_1036; // @[AesSbox.scala 40:63]
  wire  _T_1094 = _T_1038 ^ _T_1042; // @[AesSbox.scala 40:63]
  wire  _T_1096 = _T_1038 ^ _T_1064; // @[AesSbox.scala 40:63]
  wire  _T_1098 = _T_1048 ^ _T_1058; // @[AesSbox.scala 40:63]
  wire  _T_1100 = _T_1054 ^ _T_1062; // @[AesSbox.scala 40:63]
  wire  _T_1102 = _T_1056 ^ _T_1072; // @[AesSbox.scala 40:63]
  wire  _T_1104 = _T_1066 ^ _T_1078; // @[AesSbox.scala 40:63]
  wire  _T_1106 = _T_1072 ^ _T_1074; // @[AesSbox.scala 40:63]
  wire  _T_1108 = _T_1076 ^ _T_1080; // @[AesSbox.scala 40:63]
  wire  _T_1110 = _T_1072 ^ _T_1082; // @[AesSbox.scala 40:63]
  wire  _T_1112 = _T_1082 ^ _T_1084; // @[AesSbox.scala 40:63]
  wire  _T_1114 = _T_1078 ^ _T_1082; // @[AesSbox.scala 40:63]
  wire  _T_1116 = _T_1080 ^ _T_1088; // @[AesSbox.scala 40:63]
  wire  _T_1118 = _T_1086 ^ _T_1090; // @[AesSbox.scala 40:63]
  wire  _T_1120 = _T_1088 ^ _T_1104; // @[AesSbox.scala 40:63]
  wire  _T_1122 = _T_1090 ^ _T_1116; // @[AesSbox.scala 40:63]
  wire  _T_1124 = _T_1098 ^ _T_1108; // @[AesSbox.scala 40:63]
  wire  _T_1125 = _T_1094 ^ _T_1110; // @[AesSbox.scala 40:63]
  wire  _T_1126 = _T_1118 ^ _T_1124; // @[AesSbox.scala 40:63]
  wire  _T_1127 = _T_1102 ^ _T_1122; // @[AesSbox.scala 40:63]
  wire  _T_1128 = _T_1092 ^ _T_1110; // @[AesSbox.scala 40:63]
  wire  _T_1129 = _T_1112 ^ _T_1120; // @[AesSbox.scala 40:63]
  wire  _T_1130 = _T_1106 ^ _T_1114; // @[AesSbox.scala 40:63]
  wire  _T_1131 = _T_1096 ^ _T_1112; // @[AesSbox.scala 40:63]
  wire  _T_1132 = _T_1086 ^ _T_1100; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_0_3 = {_T_1125,_T_1126,_T_1127,_T_1128,_T_1129,_T_1130,_T_1131,_T_1132}; // @[Cat.scala 29:58]
  wire  _T_1158 = matrix_1_0[7] ^ matrix_1_0[4]; // @[AesSbox.scala 40:63]
  wire  _T_1160 = matrix_1_0[6] ^ matrix_1_0[4]; // @[AesSbox.scala 42:65]
  wire  _T_1161 = ~_T_1160; // @[AesSbox.scala 42:51]
  wire  _T_1163 = matrix_1_0[7] ^ matrix_1_0[6]; // @[AesSbox.scala 42:65]
  wire  _T_1164 = ~_T_1163; // @[AesSbox.scala 42:51]
  wire  _T_1166 = matrix_1_0[4] ^ matrix_1_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_1168 = matrix_1_0[3] ^ matrix_1_0[0]; // @[AesSbox.scala 42:65]
  wire  _T_1169 = ~_T_1168; // @[AesSbox.scala 42:51]
  wire  _T_1171 = matrix_1_0[1] ^ matrix_1_0[0]; // @[AesSbox.scala 40:63]
  wire  _T_1173 = matrix_1_0[6] ^ _T_1158; // @[AesSbox.scala 42:65]
  wire  _T_1174 = ~_T_1173; // @[AesSbox.scala 42:51]
  wire  _T_1176 = _T_1161 ^ _T_1171; // @[AesSbox.scala 40:63]
  wire  _T_1178 = matrix_1_0[0] ^ _T_1166; // @[AesSbox.scala 42:65]
  wire  _T_1179 = ~_T_1178; // @[AesSbox.scala 42:51]
  wire  _T_1181 = _T_1164 ^ _T_1169; // @[AesSbox.scala 40:63]
  wire  _T_1183 = _T_1164 ^ _T_1171; // @[AesSbox.scala 40:63]
  wire  _T_1185 = _T_1166 ^ _T_1171; // @[AesSbox.scala 40:63]
  wire  _T_1187 = matrix_1_0[5] ^ _T_1166; // @[AesSbox.scala 42:65]
  wire  _T_1188 = ~_T_1187; // @[AesSbox.scala 42:51]
  wire  _T_1190 = matrix_1_0[6] ^ matrix_1_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_1192 = matrix_1_0[5] ^ _T_1176; // @[AesSbox.scala 42:65]
  wire  _T_1193 = ~_T_1192; // @[AesSbox.scala 42:51]
  wire  _T_1195 = _T_1169 ^ _T_1190; // @[AesSbox.scala 40:63]
  wire  _T_1197 = matrix_1_0[3] ^ _T_1174; // @[AesSbox.scala 40:63]
  wire  _T_1199 = matrix_1_0[5] ^ matrix_1_0[2]; // @[AesSbox.scala 42:65]
  wire  _T_1200 = ~_T_1199; // @[AesSbox.scala 42:51]
  wire  _T_1202 = matrix_1_0[2] ^ matrix_1_0[1]; // @[AesSbox.scala 42:65]
  wire  _T_1203 = ~_T_1202; // @[AesSbox.scala 42:51]
  wire  _T_1205 = matrix_1_0[5] ^ matrix_1_0[3]; // @[AesSbox.scala 42:65]
  wire  _T_1206 = ~_T_1205; // @[AesSbox.scala 42:51]
  wire  _T_1208 = matrix_1_0[7] ^ _T_1200; // @[AesSbox.scala 40:63]
  wire  _T_1210 = _T_1161 ^ _T_1200; // @[AesSbox.scala 40:63]
  wire  _T_1212 = _T_1190 ^ _T_1206; // @[AesSbox.scala 40:63]
  wire  _T_1214 = _T_1166 ^ _T_1203; // @[AesSbox.scala 40:63]
  wire  _T_1216 = _T_1181 ^ _T_1214; // @[AesSbox.scala 40:63]
  wire  _T_1218 = _T_1181 ^ _T_1203; // @[AesSbox.scala 40:63]
  wire  _T_1220 = _T_1185 ^ _T_1212; // @[AesSbox.scala 40:63]
  wire  _T_1222 = _T_1183 & _T_1210; // @[AesSbox.scala 41:63]
  wire  _T_1224 = _T_1158 & _T_1174; // @[AesSbox.scala 41:63]
  wire  _T_1226 = _T_1218 ^ _T_1222; // @[AesSbox.scala 40:63]
  wire  _T_1228 = _T_1176 & _T_1208; // @[AesSbox.scala 41:63]
  wire  _T_1230 = _T_1228 ^ _T_1222; // @[AesSbox.scala 40:63]
  wire  _T_1232 = _T_1185 & _T_1212; // @[AesSbox.scala 41:63]
  wire  _T_1234 = _T_1161 & _T_1179; // @[AesSbox.scala 41:63]
  wire  _T_1236 = _T_1220 ^ _T_1232; // @[AesSbox.scala 40:63]
  wire  _T_1238 = _T_1195 & _T_1193; // @[AesSbox.scala 41:63]
  wire  _T_1240 = _T_1238 ^ _T_1232; // @[AesSbox.scala 40:63]
  wire  _T_1242 = _T_1166 & _T_1216; // @[AesSbox.scala 41:63]
  wire  _T_1244 = _T_1197 & _T_1214; // @[AesSbox.scala 41:63]
  wire  _T_1246 = _T_1244 ^ _T_1242; // @[AesSbox.scala 40:63]
  wire  _T_1248 = _T_1164 & _T_1181; // @[AesSbox.scala 41:63]
  wire  _T_1250 = _T_1248 ^ _T_1242; // @[AesSbox.scala 40:63]
  wire  _T_1252 = _T_1226 ^ _T_1224; // @[AesSbox.scala 40:63]
  wire  _T_1254 = _T_1230 ^ _T_1169; // @[AesSbox.scala 40:63]
  wire  _T_1256 = _T_1236 ^ _T_1234; // @[AesSbox.scala 40:63]
  wire  _T_1258 = _T_1240 ^ _T_1250; // @[AesSbox.scala 40:63]
  wire  _T_1260 = _T_1252 ^ _T_1246; // @[AesSbox.scala 40:63]
  wire  _T_1262 = _T_1254 ^ _T_1250; // @[AesSbox.scala 40:63]
  wire  _T_1264 = _T_1256 ^ _T_1246; // @[AesSbox.scala 40:63]
  wire  _T_1266 = _T_1258 ^ _T_1188; // @[AesSbox.scala 40:63]
  wire  _T_1268 = _T_1264 ^ _T_1266; // @[AesSbox.scala 40:63]
  wire  _T_1270 = _T_1264 & _T_1260; // @[AesSbox.scala 41:63]
  wire  _T_1272 = _T_1262 ^ _T_1270; // @[AesSbox.scala 40:63]
  wire  _T_1274 = _T_1260 ^ _T_1262; // @[AesSbox.scala 40:63]
  wire  _T_1276 = _T_1266 ^ _T_1270; // @[AesSbox.scala 40:63]
  wire  _T_1278 = _T_1276 & _T_1274; // @[AesSbox.scala 41:63]
  wire  _T_1280 = _T_1272 & _T_1268; // @[AesSbox.scala 41:63]
  wire  _T_1282 = _T_1260 & _T_1266; // @[AesSbox.scala 41:63]
  wire  _T_1284 = _T_1274 & _T_1282; // @[AesSbox.scala 41:63]
  wire  _T_1286 = _T_1274 ^ _T_1270; // @[AesSbox.scala 40:63]
  wire  _T_1288 = _T_1262 & _T_1264; // @[AesSbox.scala 41:63]
  wire  _T_1290 = _T_1268 & _T_1288; // @[AesSbox.scala 41:63]
  wire  _T_1292 = _T_1268 ^ _T_1270; // @[AesSbox.scala 40:63]
  wire  _T_1294 = _T_1262 ^ _T_1278; // @[AesSbox.scala 40:63]
  wire  _T_1296 = _T_1284 ^ _T_1286; // @[AesSbox.scala 40:63]
  wire  _T_1298 = _T_1266 ^ _T_1280; // @[AesSbox.scala 40:63]
  wire  _T_1300 = _T_1290 ^ _T_1292; // @[AesSbox.scala 40:63]
  wire  _T_1302 = _T_1296 ^ _T_1300; // @[AesSbox.scala 40:63]
  wire  _T_1304 = _T_1294 ^ _T_1298; // @[AesSbox.scala 40:63]
  wire  _T_1306 = _T_1294 ^ _T_1296; // @[AesSbox.scala 40:63]
  wire  _T_1308 = _T_1298 ^ _T_1300; // @[AesSbox.scala 40:63]
  wire  _T_1310 = _T_1304 ^ _T_1302; // @[AesSbox.scala 40:63]
  wire  _T_1312 = _T_1308 & _T_1210; // @[AesSbox.scala 41:63]
  wire  _T_1314 = _T_1300 & _T_1174; // @[AesSbox.scala 41:63]
  wire  _T_1316 = _T_1298 & _T_1208; // @[AesSbox.scala 41:63]
  wire  _T_1318 = _T_1306 & _T_1212; // @[AesSbox.scala 41:63]
  wire  _T_1320 = _T_1296 & _T_1179; // @[AesSbox.scala 41:63]
  wire  _T_1322 = _T_1294 & _T_1193; // @[AesSbox.scala 41:63]
  wire  _T_1324 = _T_1304 & _T_1216; // @[AesSbox.scala 41:63]
  wire  _T_1326 = _T_1310 & _T_1214; // @[AesSbox.scala 41:63]
  wire  _T_1328 = _T_1302 & _T_1181; // @[AesSbox.scala 41:63]
  wire  _T_1330 = _T_1308 & _T_1183; // @[AesSbox.scala 41:63]
  wire  _T_1332 = _T_1300 & _T_1158; // @[AesSbox.scala 41:63]
  wire  _T_1334 = _T_1298 & _T_1176; // @[AesSbox.scala 41:63]
  wire  _T_1336 = _T_1306 & _T_1185; // @[AesSbox.scala 41:63]
  wire  _T_1338 = _T_1296 & _T_1161; // @[AesSbox.scala 41:63]
  wire  _T_1340 = _T_1294 & _T_1195; // @[AesSbox.scala 41:63]
  wire  _T_1342 = _T_1304 & _T_1166; // @[AesSbox.scala 41:63]
  wire  _T_1344 = _T_1310 & _T_1197; // @[AesSbox.scala 41:63]
  wire  _T_1346 = _T_1302 & _T_1164; // @[AesSbox.scala 41:63]
  wire  _T_1348 = _T_1324 ^ _T_1342; // @[AesSbox.scala 40:63]
  wire  _T_1350 = _T_1336 ^ _T_1338; // @[AesSbox.scala 40:63]
  wire  _T_1352 = _T_1328 ^ _T_1344; // @[AesSbox.scala 40:63]
  wire  _T_1354 = _T_1314 ^ _T_1320; // @[AesSbox.scala 40:63]
  wire  _T_1356 = _T_1316 ^ _T_1332; // @[AesSbox.scala 40:63]
  wire  _T_1358 = _T_1312 ^ _T_1322; // @[AesSbox.scala 40:63]
  wire  _T_1360 = _T_1318 ^ _T_1340; // @[AesSbox.scala 40:63]
  wire  _T_1362 = _T_1348 ^ _T_1350; // @[AesSbox.scala 40:63]
  wire  _T_1364 = _T_1320 ^ _T_1326; // @[AesSbox.scala 40:63]
  wire  _T_1366 = _T_1330 ^ _T_1346; // @[AesSbox.scala 40:63]
  wire  _T_1368 = _T_1334 ^ _T_1356; // @[AesSbox.scala 40:63]
  wire  _T_1370 = _T_1348 ^ _T_1354; // @[AesSbox.scala 40:63]
  wire  _T_1372 = _T_1312 ^ _T_1316; // @[AesSbox.scala 40:63]
  wire  _T_1374 = _T_1318 ^ _T_1322; // @[AesSbox.scala 40:63]
  wire  _T_1376 = _T_1318 ^ _T_1344; // @[AesSbox.scala 40:63]
  wire  _T_1378 = _T_1328 ^ _T_1338; // @[AesSbox.scala 40:63]
  wire  _T_1380 = _T_1334 ^ _T_1342; // @[AesSbox.scala 40:63]
  wire  _T_1382 = _T_1336 ^ _T_1352; // @[AesSbox.scala 40:63]
  wire  _T_1384 = _T_1346 ^ _T_1358; // @[AesSbox.scala 40:63]
  wire  _T_1386 = _T_1352 ^ _T_1354; // @[AesSbox.scala 40:63]
  wire  _T_1388 = _T_1356 ^ _T_1360; // @[AesSbox.scala 40:63]
  wire  _T_1390 = _T_1352 ^ _T_1362; // @[AesSbox.scala 40:63]
  wire  _T_1392 = _T_1362 ^ _T_1364; // @[AesSbox.scala 40:63]
  wire  _T_1394 = _T_1358 ^ _T_1362; // @[AesSbox.scala 40:63]
  wire  _T_1396 = _T_1360 ^ _T_1368; // @[AesSbox.scala 40:63]
  wire  _T_1398 = _T_1366 ^ _T_1370; // @[AesSbox.scala 40:63]
  wire  _T_1400 = _T_1368 ^ _T_1384; // @[AesSbox.scala 40:63]
  wire  _T_1402 = _T_1370 ^ _T_1396; // @[AesSbox.scala 40:63]
  wire  _T_1404 = _T_1378 ^ _T_1388; // @[AesSbox.scala 40:63]
  wire  _T_1405 = _T_1374 ^ _T_1390; // @[AesSbox.scala 40:63]
  wire  _T_1406 = _T_1398 ^ _T_1404; // @[AesSbox.scala 40:63]
  wire  _T_1407 = _T_1382 ^ _T_1402; // @[AesSbox.scala 40:63]
  wire  _T_1408 = _T_1372 ^ _T_1390; // @[AesSbox.scala 40:63]
  wire  _T_1409 = _T_1392 ^ _T_1400; // @[AesSbox.scala 40:63]
  wire  _T_1410 = _T_1386 ^ _T_1394; // @[AesSbox.scala 40:63]
  wire  _T_1411 = _T_1376 ^ _T_1392; // @[AesSbox.scala 40:63]
  wire  _T_1412 = _T_1366 ^ _T_1380; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_1_0 = {_T_1405,_T_1406,_T_1407,_T_1408,_T_1409,_T_1410,_T_1411,_T_1412}; // @[Cat.scala 29:58]
  wire  _T_1437 = matrix_0_1[7] ^ matrix_0_1[4]; // @[AesSbox.scala 40:63]
  wire  _T_1439 = matrix_0_1[6] ^ matrix_0_1[4]; // @[AesSbox.scala 42:65]
  wire  _T_1440 = ~_T_1439; // @[AesSbox.scala 42:51]
  wire  _T_1442 = matrix_0_1[7] ^ matrix_0_1[6]; // @[AesSbox.scala 42:65]
  wire  _T_1443 = ~_T_1442; // @[AesSbox.scala 42:51]
  wire  _T_1445 = matrix_0_1[4] ^ matrix_0_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_1447 = matrix_0_1[3] ^ matrix_0_1[0]; // @[AesSbox.scala 42:65]
  wire  _T_1448 = ~_T_1447; // @[AesSbox.scala 42:51]
  wire  _T_1450 = matrix_0_1[1] ^ matrix_0_1[0]; // @[AesSbox.scala 40:63]
  wire  _T_1452 = matrix_0_1[6] ^ _T_1437; // @[AesSbox.scala 42:65]
  wire  _T_1453 = ~_T_1452; // @[AesSbox.scala 42:51]
  wire  _T_1455 = _T_1440 ^ _T_1450; // @[AesSbox.scala 40:63]
  wire  _T_1457 = matrix_0_1[0] ^ _T_1445; // @[AesSbox.scala 42:65]
  wire  _T_1458 = ~_T_1457; // @[AesSbox.scala 42:51]
  wire  _T_1460 = _T_1443 ^ _T_1448; // @[AesSbox.scala 40:63]
  wire  _T_1462 = _T_1443 ^ _T_1450; // @[AesSbox.scala 40:63]
  wire  _T_1464 = _T_1445 ^ _T_1450; // @[AesSbox.scala 40:63]
  wire  _T_1466 = matrix_0_1[5] ^ _T_1445; // @[AesSbox.scala 42:65]
  wire  _T_1467 = ~_T_1466; // @[AesSbox.scala 42:51]
  wire  _T_1469 = matrix_0_1[6] ^ matrix_0_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_1471 = matrix_0_1[5] ^ _T_1455; // @[AesSbox.scala 42:65]
  wire  _T_1472 = ~_T_1471; // @[AesSbox.scala 42:51]
  wire  _T_1474 = _T_1448 ^ _T_1469; // @[AesSbox.scala 40:63]
  wire  _T_1476 = matrix_0_1[3] ^ _T_1453; // @[AesSbox.scala 40:63]
  wire  _T_1478 = matrix_0_1[5] ^ matrix_0_1[2]; // @[AesSbox.scala 42:65]
  wire  _T_1479 = ~_T_1478; // @[AesSbox.scala 42:51]
  wire  _T_1481 = matrix_0_1[2] ^ matrix_0_1[1]; // @[AesSbox.scala 42:65]
  wire  _T_1482 = ~_T_1481; // @[AesSbox.scala 42:51]
  wire  _T_1484 = matrix_0_1[5] ^ matrix_0_1[3]; // @[AesSbox.scala 42:65]
  wire  _T_1485 = ~_T_1484; // @[AesSbox.scala 42:51]
  wire  _T_1487 = matrix_0_1[7] ^ _T_1479; // @[AesSbox.scala 40:63]
  wire  _T_1489 = _T_1440 ^ _T_1479; // @[AesSbox.scala 40:63]
  wire  _T_1491 = _T_1469 ^ _T_1485; // @[AesSbox.scala 40:63]
  wire  _T_1493 = _T_1445 ^ _T_1482; // @[AesSbox.scala 40:63]
  wire  _T_1495 = _T_1460 ^ _T_1493; // @[AesSbox.scala 40:63]
  wire  _T_1497 = _T_1460 ^ _T_1482; // @[AesSbox.scala 40:63]
  wire  _T_1499 = _T_1464 ^ _T_1491; // @[AesSbox.scala 40:63]
  wire  _T_1501 = _T_1462 & _T_1489; // @[AesSbox.scala 41:63]
  wire  _T_1503 = _T_1437 & _T_1453; // @[AesSbox.scala 41:63]
  wire  _T_1505 = _T_1497 ^ _T_1501; // @[AesSbox.scala 40:63]
  wire  _T_1507 = _T_1455 & _T_1487; // @[AesSbox.scala 41:63]
  wire  _T_1509 = _T_1507 ^ _T_1501; // @[AesSbox.scala 40:63]
  wire  _T_1511 = _T_1464 & _T_1491; // @[AesSbox.scala 41:63]
  wire  _T_1513 = _T_1440 & _T_1458; // @[AesSbox.scala 41:63]
  wire  _T_1515 = _T_1499 ^ _T_1511; // @[AesSbox.scala 40:63]
  wire  _T_1517 = _T_1474 & _T_1472; // @[AesSbox.scala 41:63]
  wire  _T_1519 = _T_1517 ^ _T_1511; // @[AesSbox.scala 40:63]
  wire  _T_1521 = _T_1445 & _T_1495; // @[AesSbox.scala 41:63]
  wire  _T_1523 = _T_1476 & _T_1493; // @[AesSbox.scala 41:63]
  wire  _T_1525 = _T_1523 ^ _T_1521; // @[AesSbox.scala 40:63]
  wire  _T_1527 = _T_1443 & _T_1460; // @[AesSbox.scala 41:63]
  wire  _T_1529 = _T_1527 ^ _T_1521; // @[AesSbox.scala 40:63]
  wire  _T_1531 = _T_1505 ^ _T_1503; // @[AesSbox.scala 40:63]
  wire  _T_1533 = _T_1509 ^ _T_1448; // @[AesSbox.scala 40:63]
  wire  _T_1535 = _T_1515 ^ _T_1513; // @[AesSbox.scala 40:63]
  wire  _T_1537 = _T_1519 ^ _T_1529; // @[AesSbox.scala 40:63]
  wire  _T_1539 = _T_1531 ^ _T_1525; // @[AesSbox.scala 40:63]
  wire  _T_1541 = _T_1533 ^ _T_1529; // @[AesSbox.scala 40:63]
  wire  _T_1543 = _T_1535 ^ _T_1525; // @[AesSbox.scala 40:63]
  wire  _T_1545 = _T_1537 ^ _T_1467; // @[AesSbox.scala 40:63]
  wire  _T_1547 = _T_1543 ^ _T_1545; // @[AesSbox.scala 40:63]
  wire  _T_1549 = _T_1543 & _T_1539; // @[AesSbox.scala 41:63]
  wire  _T_1551 = _T_1541 ^ _T_1549; // @[AesSbox.scala 40:63]
  wire  _T_1553 = _T_1539 ^ _T_1541; // @[AesSbox.scala 40:63]
  wire  _T_1555 = _T_1545 ^ _T_1549; // @[AesSbox.scala 40:63]
  wire  _T_1557 = _T_1555 & _T_1553; // @[AesSbox.scala 41:63]
  wire  _T_1559 = _T_1551 & _T_1547; // @[AesSbox.scala 41:63]
  wire  _T_1561 = _T_1539 & _T_1545; // @[AesSbox.scala 41:63]
  wire  _T_1563 = _T_1553 & _T_1561; // @[AesSbox.scala 41:63]
  wire  _T_1565 = _T_1553 ^ _T_1549; // @[AesSbox.scala 40:63]
  wire  _T_1567 = _T_1541 & _T_1543; // @[AesSbox.scala 41:63]
  wire  _T_1569 = _T_1547 & _T_1567; // @[AesSbox.scala 41:63]
  wire  _T_1571 = _T_1547 ^ _T_1549; // @[AesSbox.scala 40:63]
  wire  _T_1573 = _T_1541 ^ _T_1557; // @[AesSbox.scala 40:63]
  wire  _T_1575 = _T_1563 ^ _T_1565; // @[AesSbox.scala 40:63]
  wire  _T_1577 = _T_1545 ^ _T_1559; // @[AesSbox.scala 40:63]
  wire  _T_1579 = _T_1569 ^ _T_1571; // @[AesSbox.scala 40:63]
  wire  _T_1581 = _T_1575 ^ _T_1579; // @[AesSbox.scala 40:63]
  wire  _T_1583 = _T_1573 ^ _T_1577; // @[AesSbox.scala 40:63]
  wire  _T_1585 = _T_1573 ^ _T_1575; // @[AesSbox.scala 40:63]
  wire  _T_1587 = _T_1577 ^ _T_1579; // @[AesSbox.scala 40:63]
  wire  _T_1589 = _T_1583 ^ _T_1581; // @[AesSbox.scala 40:63]
  wire  _T_1591 = _T_1587 & _T_1489; // @[AesSbox.scala 41:63]
  wire  _T_1593 = _T_1579 & _T_1453; // @[AesSbox.scala 41:63]
  wire  _T_1595 = _T_1577 & _T_1487; // @[AesSbox.scala 41:63]
  wire  _T_1597 = _T_1585 & _T_1491; // @[AesSbox.scala 41:63]
  wire  _T_1599 = _T_1575 & _T_1458; // @[AesSbox.scala 41:63]
  wire  _T_1601 = _T_1573 & _T_1472; // @[AesSbox.scala 41:63]
  wire  _T_1603 = _T_1583 & _T_1495; // @[AesSbox.scala 41:63]
  wire  _T_1605 = _T_1589 & _T_1493; // @[AesSbox.scala 41:63]
  wire  _T_1607 = _T_1581 & _T_1460; // @[AesSbox.scala 41:63]
  wire  _T_1609 = _T_1587 & _T_1462; // @[AesSbox.scala 41:63]
  wire  _T_1611 = _T_1579 & _T_1437; // @[AesSbox.scala 41:63]
  wire  _T_1613 = _T_1577 & _T_1455; // @[AesSbox.scala 41:63]
  wire  _T_1615 = _T_1585 & _T_1464; // @[AesSbox.scala 41:63]
  wire  _T_1617 = _T_1575 & _T_1440; // @[AesSbox.scala 41:63]
  wire  _T_1619 = _T_1573 & _T_1474; // @[AesSbox.scala 41:63]
  wire  _T_1621 = _T_1583 & _T_1445; // @[AesSbox.scala 41:63]
  wire  _T_1623 = _T_1589 & _T_1476; // @[AesSbox.scala 41:63]
  wire  _T_1625 = _T_1581 & _T_1443; // @[AesSbox.scala 41:63]
  wire  _T_1627 = _T_1603 ^ _T_1621; // @[AesSbox.scala 40:63]
  wire  _T_1629 = _T_1615 ^ _T_1617; // @[AesSbox.scala 40:63]
  wire  _T_1631 = _T_1607 ^ _T_1623; // @[AesSbox.scala 40:63]
  wire  _T_1633 = _T_1593 ^ _T_1599; // @[AesSbox.scala 40:63]
  wire  _T_1635 = _T_1595 ^ _T_1611; // @[AesSbox.scala 40:63]
  wire  _T_1637 = _T_1591 ^ _T_1601; // @[AesSbox.scala 40:63]
  wire  _T_1639 = _T_1597 ^ _T_1619; // @[AesSbox.scala 40:63]
  wire  _T_1641 = _T_1627 ^ _T_1629; // @[AesSbox.scala 40:63]
  wire  _T_1643 = _T_1599 ^ _T_1605; // @[AesSbox.scala 40:63]
  wire  _T_1645 = _T_1609 ^ _T_1625; // @[AesSbox.scala 40:63]
  wire  _T_1647 = _T_1613 ^ _T_1635; // @[AesSbox.scala 40:63]
  wire  _T_1649 = _T_1627 ^ _T_1633; // @[AesSbox.scala 40:63]
  wire  _T_1651 = _T_1591 ^ _T_1595; // @[AesSbox.scala 40:63]
  wire  _T_1653 = _T_1597 ^ _T_1601; // @[AesSbox.scala 40:63]
  wire  _T_1655 = _T_1597 ^ _T_1623; // @[AesSbox.scala 40:63]
  wire  _T_1657 = _T_1607 ^ _T_1617; // @[AesSbox.scala 40:63]
  wire  _T_1659 = _T_1613 ^ _T_1621; // @[AesSbox.scala 40:63]
  wire  _T_1661 = _T_1615 ^ _T_1631; // @[AesSbox.scala 40:63]
  wire  _T_1663 = _T_1625 ^ _T_1637; // @[AesSbox.scala 40:63]
  wire  _T_1665 = _T_1631 ^ _T_1633; // @[AesSbox.scala 40:63]
  wire  _T_1667 = _T_1635 ^ _T_1639; // @[AesSbox.scala 40:63]
  wire  _T_1669 = _T_1631 ^ _T_1641; // @[AesSbox.scala 40:63]
  wire  _T_1671 = _T_1641 ^ _T_1643; // @[AesSbox.scala 40:63]
  wire  _T_1673 = _T_1637 ^ _T_1641; // @[AesSbox.scala 40:63]
  wire  _T_1675 = _T_1639 ^ _T_1647; // @[AesSbox.scala 40:63]
  wire  _T_1677 = _T_1645 ^ _T_1649; // @[AesSbox.scala 40:63]
  wire  _T_1679 = _T_1647 ^ _T_1663; // @[AesSbox.scala 40:63]
  wire  _T_1681 = _T_1649 ^ _T_1675; // @[AesSbox.scala 40:63]
  wire  _T_1683 = _T_1657 ^ _T_1667; // @[AesSbox.scala 40:63]
  wire  _T_1684 = _T_1653 ^ _T_1669; // @[AesSbox.scala 40:63]
  wire  _T_1685 = _T_1677 ^ _T_1683; // @[AesSbox.scala 40:63]
  wire  _T_1686 = _T_1661 ^ _T_1681; // @[AesSbox.scala 40:63]
  wire  _T_1687 = _T_1651 ^ _T_1669; // @[AesSbox.scala 40:63]
  wire  _T_1688 = _T_1671 ^ _T_1679; // @[AesSbox.scala 40:63]
  wire  _T_1689 = _T_1665 ^ _T_1673; // @[AesSbox.scala 40:63]
  wire  _T_1690 = _T_1655 ^ _T_1671; // @[AesSbox.scala 40:63]
  wire  _T_1691 = _T_1645 ^ _T_1659; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_1_1 = {_T_1684,_T_1685,_T_1686,_T_1687,_T_1688,_T_1689,_T_1690,_T_1691}; // @[Cat.scala 29:58]
  wire  _T_1716 = matrix_3_2[7] ^ matrix_3_2[4]; // @[AesSbox.scala 40:63]
  wire  _T_1718 = matrix_3_2[6] ^ matrix_3_2[4]; // @[AesSbox.scala 42:65]
  wire  _T_1719 = ~_T_1718; // @[AesSbox.scala 42:51]
  wire  _T_1721 = matrix_3_2[7] ^ matrix_3_2[6]; // @[AesSbox.scala 42:65]
  wire  _T_1722 = ~_T_1721; // @[AesSbox.scala 42:51]
  wire  _T_1724 = matrix_3_2[4] ^ matrix_3_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_1726 = matrix_3_2[3] ^ matrix_3_2[0]; // @[AesSbox.scala 42:65]
  wire  _T_1727 = ~_T_1726; // @[AesSbox.scala 42:51]
  wire  _T_1729 = matrix_3_2[1] ^ matrix_3_2[0]; // @[AesSbox.scala 40:63]
  wire  _T_1731 = matrix_3_2[6] ^ _T_1716; // @[AesSbox.scala 42:65]
  wire  _T_1732 = ~_T_1731; // @[AesSbox.scala 42:51]
  wire  _T_1734 = _T_1719 ^ _T_1729; // @[AesSbox.scala 40:63]
  wire  _T_1736 = matrix_3_2[0] ^ _T_1724; // @[AesSbox.scala 42:65]
  wire  _T_1737 = ~_T_1736; // @[AesSbox.scala 42:51]
  wire  _T_1739 = _T_1722 ^ _T_1727; // @[AesSbox.scala 40:63]
  wire  _T_1741 = _T_1722 ^ _T_1729; // @[AesSbox.scala 40:63]
  wire  _T_1743 = _T_1724 ^ _T_1729; // @[AesSbox.scala 40:63]
  wire  _T_1745 = matrix_3_2[5] ^ _T_1724; // @[AesSbox.scala 42:65]
  wire  _T_1746 = ~_T_1745; // @[AesSbox.scala 42:51]
  wire  _T_1748 = matrix_3_2[6] ^ matrix_3_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_1750 = matrix_3_2[5] ^ _T_1734; // @[AesSbox.scala 42:65]
  wire  _T_1751 = ~_T_1750; // @[AesSbox.scala 42:51]
  wire  _T_1753 = _T_1727 ^ _T_1748; // @[AesSbox.scala 40:63]
  wire  _T_1755 = matrix_3_2[3] ^ _T_1732; // @[AesSbox.scala 40:63]
  wire  _T_1757 = matrix_3_2[5] ^ matrix_3_2[2]; // @[AesSbox.scala 42:65]
  wire  _T_1758 = ~_T_1757; // @[AesSbox.scala 42:51]
  wire  _T_1760 = matrix_3_2[2] ^ matrix_3_2[1]; // @[AesSbox.scala 42:65]
  wire  _T_1761 = ~_T_1760; // @[AesSbox.scala 42:51]
  wire  _T_1763 = matrix_3_2[5] ^ matrix_3_2[3]; // @[AesSbox.scala 42:65]
  wire  _T_1764 = ~_T_1763; // @[AesSbox.scala 42:51]
  wire  _T_1766 = matrix_3_2[7] ^ _T_1758; // @[AesSbox.scala 40:63]
  wire  _T_1768 = _T_1719 ^ _T_1758; // @[AesSbox.scala 40:63]
  wire  _T_1770 = _T_1748 ^ _T_1764; // @[AesSbox.scala 40:63]
  wire  _T_1772 = _T_1724 ^ _T_1761; // @[AesSbox.scala 40:63]
  wire  _T_1774 = _T_1739 ^ _T_1772; // @[AesSbox.scala 40:63]
  wire  _T_1776 = _T_1739 ^ _T_1761; // @[AesSbox.scala 40:63]
  wire  _T_1778 = _T_1743 ^ _T_1770; // @[AesSbox.scala 40:63]
  wire  _T_1780 = _T_1741 & _T_1768; // @[AesSbox.scala 41:63]
  wire  _T_1782 = _T_1716 & _T_1732; // @[AesSbox.scala 41:63]
  wire  _T_1784 = _T_1776 ^ _T_1780; // @[AesSbox.scala 40:63]
  wire  _T_1786 = _T_1734 & _T_1766; // @[AesSbox.scala 41:63]
  wire  _T_1788 = _T_1786 ^ _T_1780; // @[AesSbox.scala 40:63]
  wire  _T_1790 = _T_1743 & _T_1770; // @[AesSbox.scala 41:63]
  wire  _T_1792 = _T_1719 & _T_1737; // @[AesSbox.scala 41:63]
  wire  _T_1794 = _T_1778 ^ _T_1790; // @[AesSbox.scala 40:63]
  wire  _T_1796 = _T_1753 & _T_1751; // @[AesSbox.scala 41:63]
  wire  _T_1798 = _T_1796 ^ _T_1790; // @[AesSbox.scala 40:63]
  wire  _T_1800 = _T_1724 & _T_1774; // @[AesSbox.scala 41:63]
  wire  _T_1802 = _T_1755 & _T_1772; // @[AesSbox.scala 41:63]
  wire  _T_1804 = _T_1802 ^ _T_1800; // @[AesSbox.scala 40:63]
  wire  _T_1806 = _T_1722 & _T_1739; // @[AesSbox.scala 41:63]
  wire  _T_1808 = _T_1806 ^ _T_1800; // @[AesSbox.scala 40:63]
  wire  _T_1810 = _T_1784 ^ _T_1782; // @[AesSbox.scala 40:63]
  wire  _T_1812 = _T_1788 ^ _T_1727; // @[AesSbox.scala 40:63]
  wire  _T_1814 = _T_1794 ^ _T_1792; // @[AesSbox.scala 40:63]
  wire  _T_1816 = _T_1798 ^ _T_1808; // @[AesSbox.scala 40:63]
  wire  _T_1818 = _T_1810 ^ _T_1804; // @[AesSbox.scala 40:63]
  wire  _T_1820 = _T_1812 ^ _T_1808; // @[AesSbox.scala 40:63]
  wire  _T_1822 = _T_1814 ^ _T_1804; // @[AesSbox.scala 40:63]
  wire  _T_1824 = _T_1816 ^ _T_1746; // @[AesSbox.scala 40:63]
  wire  _T_1826 = _T_1822 ^ _T_1824; // @[AesSbox.scala 40:63]
  wire  _T_1828 = _T_1822 & _T_1818; // @[AesSbox.scala 41:63]
  wire  _T_1830 = _T_1820 ^ _T_1828; // @[AesSbox.scala 40:63]
  wire  _T_1832 = _T_1818 ^ _T_1820; // @[AesSbox.scala 40:63]
  wire  _T_1834 = _T_1824 ^ _T_1828; // @[AesSbox.scala 40:63]
  wire  _T_1836 = _T_1834 & _T_1832; // @[AesSbox.scala 41:63]
  wire  _T_1838 = _T_1830 & _T_1826; // @[AesSbox.scala 41:63]
  wire  _T_1840 = _T_1818 & _T_1824; // @[AesSbox.scala 41:63]
  wire  _T_1842 = _T_1832 & _T_1840; // @[AesSbox.scala 41:63]
  wire  _T_1844 = _T_1832 ^ _T_1828; // @[AesSbox.scala 40:63]
  wire  _T_1846 = _T_1820 & _T_1822; // @[AesSbox.scala 41:63]
  wire  _T_1848 = _T_1826 & _T_1846; // @[AesSbox.scala 41:63]
  wire  _T_1850 = _T_1826 ^ _T_1828; // @[AesSbox.scala 40:63]
  wire  _T_1852 = _T_1820 ^ _T_1836; // @[AesSbox.scala 40:63]
  wire  _T_1854 = _T_1842 ^ _T_1844; // @[AesSbox.scala 40:63]
  wire  _T_1856 = _T_1824 ^ _T_1838; // @[AesSbox.scala 40:63]
  wire  _T_1858 = _T_1848 ^ _T_1850; // @[AesSbox.scala 40:63]
  wire  _T_1860 = _T_1854 ^ _T_1858; // @[AesSbox.scala 40:63]
  wire  _T_1862 = _T_1852 ^ _T_1856; // @[AesSbox.scala 40:63]
  wire  _T_1864 = _T_1852 ^ _T_1854; // @[AesSbox.scala 40:63]
  wire  _T_1866 = _T_1856 ^ _T_1858; // @[AesSbox.scala 40:63]
  wire  _T_1868 = _T_1862 ^ _T_1860; // @[AesSbox.scala 40:63]
  wire  _T_1870 = _T_1866 & _T_1768; // @[AesSbox.scala 41:63]
  wire  _T_1872 = _T_1858 & _T_1732; // @[AesSbox.scala 41:63]
  wire  _T_1874 = _T_1856 & _T_1766; // @[AesSbox.scala 41:63]
  wire  _T_1876 = _T_1864 & _T_1770; // @[AesSbox.scala 41:63]
  wire  _T_1878 = _T_1854 & _T_1737; // @[AesSbox.scala 41:63]
  wire  _T_1880 = _T_1852 & _T_1751; // @[AesSbox.scala 41:63]
  wire  _T_1882 = _T_1862 & _T_1774; // @[AesSbox.scala 41:63]
  wire  _T_1884 = _T_1868 & _T_1772; // @[AesSbox.scala 41:63]
  wire  _T_1886 = _T_1860 & _T_1739; // @[AesSbox.scala 41:63]
  wire  _T_1888 = _T_1866 & _T_1741; // @[AesSbox.scala 41:63]
  wire  _T_1890 = _T_1858 & _T_1716; // @[AesSbox.scala 41:63]
  wire  _T_1892 = _T_1856 & _T_1734; // @[AesSbox.scala 41:63]
  wire  _T_1894 = _T_1864 & _T_1743; // @[AesSbox.scala 41:63]
  wire  _T_1896 = _T_1854 & _T_1719; // @[AesSbox.scala 41:63]
  wire  _T_1898 = _T_1852 & _T_1753; // @[AesSbox.scala 41:63]
  wire  _T_1900 = _T_1862 & _T_1724; // @[AesSbox.scala 41:63]
  wire  _T_1902 = _T_1868 & _T_1755; // @[AesSbox.scala 41:63]
  wire  _T_1904 = _T_1860 & _T_1722; // @[AesSbox.scala 41:63]
  wire  _T_1906 = _T_1882 ^ _T_1900; // @[AesSbox.scala 40:63]
  wire  _T_1908 = _T_1894 ^ _T_1896; // @[AesSbox.scala 40:63]
  wire  _T_1910 = _T_1886 ^ _T_1902; // @[AesSbox.scala 40:63]
  wire  _T_1912 = _T_1872 ^ _T_1878; // @[AesSbox.scala 40:63]
  wire  _T_1914 = _T_1874 ^ _T_1890; // @[AesSbox.scala 40:63]
  wire  _T_1916 = _T_1870 ^ _T_1880; // @[AesSbox.scala 40:63]
  wire  _T_1918 = _T_1876 ^ _T_1898; // @[AesSbox.scala 40:63]
  wire  _T_1920 = _T_1906 ^ _T_1908; // @[AesSbox.scala 40:63]
  wire  _T_1922 = _T_1878 ^ _T_1884; // @[AesSbox.scala 40:63]
  wire  _T_1924 = _T_1888 ^ _T_1904; // @[AesSbox.scala 40:63]
  wire  _T_1926 = _T_1892 ^ _T_1914; // @[AesSbox.scala 40:63]
  wire  _T_1928 = _T_1906 ^ _T_1912; // @[AesSbox.scala 40:63]
  wire  _T_1930 = _T_1870 ^ _T_1874; // @[AesSbox.scala 40:63]
  wire  _T_1932 = _T_1876 ^ _T_1880; // @[AesSbox.scala 40:63]
  wire  _T_1934 = _T_1876 ^ _T_1902; // @[AesSbox.scala 40:63]
  wire  _T_1936 = _T_1886 ^ _T_1896; // @[AesSbox.scala 40:63]
  wire  _T_1938 = _T_1892 ^ _T_1900; // @[AesSbox.scala 40:63]
  wire  _T_1940 = _T_1894 ^ _T_1910; // @[AesSbox.scala 40:63]
  wire  _T_1942 = _T_1904 ^ _T_1916; // @[AesSbox.scala 40:63]
  wire  _T_1944 = _T_1910 ^ _T_1912; // @[AesSbox.scala 40:63]
  wire  _T_1946 = _T_1914 ^ _T_1918; // @[AesSbox.scala 40:63]
  wire  _T_1948 = _T_1910 ^ _T_1920; // @[AesSbox.scala 40:63]
  wire  _T_1950 = _T_1920 ^ _T_1922; // @[AesSbox.scala 40:63]
  wire  _T_1952 = _T_1916 ^ _T_1920; // @[AesSbox.scala 40:63]
  wire  _T_1954 = _T_1918 ^ _T_1926; // @[AesSbox.scala 40:63]
  wire  _T_1956 = _T_1924 ^ _T_1928; // @[AesSbox.scala 40:63]
  wire  _T_1958 = _T_1926 ^ _T_1942; // @[AesSbox.scala 40:63]
  wire  _T_1960 = _T_1928 ^ _T_1954; // @[AesSbox.scala 40:63]
  wire  _T_1962 = _T_1936 ^ _T_1946; // @[AesSbox.scala 40:63]
  wire  _T_1963 = _T_1932 ^ _T_1948; // @[AesSbox.scala 40:63]
  wire  _T_1964 = _T_1956 ^ _T_1962; // @[AesSbox.scala 40:63]
  wire  _T_1965 = _T_1940 ^ _T_1960; // @[AesSbox.scala 40:63]
  wire  _T_1966 = _T_1930 ^ _T_1948; // @[AesSbox.scala 40:63]
  wire  _T_1967 = _T_1950 ^ _T_1958; // @[AesSbox.scala 40:63]
  wire  _T_1968 = _T_1944 ^ _T_1952; // @[AesSbox.scala 40:63]
  wire  _T_1969 = _T_1934 ^ _T_1950; // @[AesSbox.scala 40:63]
  wire  _T_1970 = _T_1924 ^ _T_1938; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_1_2 = {_T_1963,_T_1964,_T_1965,_T_1966,_T_1967,_T_1968,_T_1969,_T_1970}; // @[Cat.scala 29:58]
  wire  _T_1995 = matrix_2_3[7] ^ matrix_2_3[4]; // @[AesSbox.scala 40:63]
  wire  _T_1997 = matrix_2_3[6] ^ matrix_2_3[4]; // @[AesSbox.scala 42:65]
  wire  _T_1998 = ~_T_1997; // @[AesSbox.scala 42:51]
  wire  _T_2000 = matrix_2_3[7] ^ matrix_2_3[6]; // @[AesSbox.scala 42:65]
  wire  _T_2001 = ~_T_2000; // @[AesSbox.scala 42:51]
  wire  _T_2003 = matrix_2_3[4] ^ matrix_2_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_2005 = matrix_2_3[3] ^ matrix_2_3[0]; // @[AesSbox.scala 42:65]
  wire  _T_2006 = ~_T_2005; // @[AesSbox.scala 42:51]
  wire  _T_2008 = matrix_2_3[1] ^ matrix_2_3[0]; // @[AesSbox.scala 40:63]
  wire  _T_2010 = matrix_2_3[6] ^ _T_1995; // @[AesSbox.scala 42:65]
  wire  _T_2011 = ~_T_2010; // @[AesSbox.scala 42:51]
  wire  _T_2013 = _T_1998 ^ _T_2008; // @[AesSbox.scala 40:63]
  wire  _T_2015 = matrix_2_3[0] ^ _T_2003; // @[AesSbox.scala 42:65]
  wire  _T_2016 = ~_T_2015; // @[AesSbox.scala 42:51]
  wire  _T_2018 = _T_2001 ^ _T_2006; // @[AesSbox.scala 40:63]
  wire  _T_2020 = _T_2001 ^ _T_2008; // @[AesSbox.scala 40:63]
  wire  _T_2022 = _T_2003 ^ _T_2008; // @[AesSbox.scala 40:63]
  wire  _T_2024 = matrix_2_3[5] ^ _T_2003; // @[AesSbox.scala 42:65]
  wire  _T_2025 = ~_T_2024; // @[AesSbox.scala 42:51]
  wire  _T_2027 = matrix_2_3[6] ^ matrix_2_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_2029 = matrix_2_3[5] ^ _T_2013; // @[AesSbox.scala 42:65]
  wire  _T_2030 = ~_T_2029; // @[AesSbox.scala 42:51]
  wire  _T_2032 = _T_2006 ^ _T_2027; // @[AesSbox.scala 40:63]
  wire  _T_2034 = matrix_2_3[3] ^ _T_2011; // @[AesSbox.scala 40:63]
  wire  _T_2036 = matrix_2_3[5] ^ matrix_2_3[2]; // @[AesSbox.scala 42:65]
  wire  _T_2037 = ~_T_2036; // @[AesSbox.scala 42:51]
  wire  _T_2039 = matrix_2_3[2] ^ matrix_2_3[1]; // @[AesSbox.scala 42:65]
  wire  _T_2040 = ~_T_2039; // @[AesSbox.scala 42:51]
  wire  _T_2042 = matrix_2_3[5] ^ matrix_2_3[3]; // @[AesSbox.scala 42:65]
  wire  _T_2043 = ~_T_2042; // @[AesSbox.scala 42:51]
  wire  _T_2045 = matrix_2_3[7] ^ _T_2037; // @[AesSbox.scala 40:63]
  wire  _T_2047 = _T_1998 ^ _T_2037; // @[AesSbox.scala 40:63]
  wire  _T_2049 = _T_2027 ^ _T_2043; // @[AesSbox.scala 40:63]
  wire  _T_2051 = _T_2003 ^ _T_2040; // @[AesSbox.scala 40:63]
  wire  _T_2053 = _T_2018 ^ _T_2051; // @[AesSbox.scala 40:63]
  wire  _T_2055 = _T_2018 ^ _T_2040; // @[AesSbox.scala 40:63]
  wire  _T_2057 = _T_2022 ^ _T_2049; // @[AesSbox.scala 40:63]
  wire  _T_2059 = _T_2020 & _T_2047; // @[AesSbox.scala 41:63]
  wire  _T_2061 = _T_1995 & _T_2011; // @[AesSbox.scala 41:63]
  wire  _T_2063 = _T_2055 ^ _T_2059; // @[AesSbox.scala 40:63]
  wire  _T_2065 = _T_2013 & _T_2045; // @[AesSbox.scala 41:63]
  wire  _T_2067 = _T_2065 ^ _T_2059; // @[AesSbox.scala 40:63]
  wire  _T_2069 = _T_2022 & _T_2049; // @[AesSbox.scala 41:63]
  wire  _T_2071 = _T_1998 & _T_2016; // @[AesSbox.scala 41:63]
  wire  _T_2073 = _T_2057 ^ _T_2069; // @[AesSbox.scala 40:63]
  wire  _T_2075 = _T_2032 & _T_2030; // @[AesSbox.scala 41:63]
  wire  _T_2077 = _T_2075 ^ _T_2069; // @[AesSbox.scala 40:63]
  wire  _T_2079 = _T_2003 & _T_2053; // @[AesSbox.scala 41:63]
  wire  _T_2081 = _T_2034 & _T_2051; // @[AesSbox.scala 41:63]
  wire  _T_2083 = _T_2081 ^ _T_2079; // @[AesSbox.scala 40:63]
  wire  _T_2085 = _T_2001 & _T_2018; // @[AesSbox.scala 41:63]
  wire  _T_2087 = _T_2085 ^ _T_2079; // @[AesSbox.scala 40:63]
  wire  _T_2089 = _T_2063 ^ _T_2061; // @[AesSbox.scala 40:63]
  wire  _T_2091 = _T_2067 ^ _T_2006; // @[AesSbox.scala 40:63]
  wire  _T_2093 = _T_2073 ^ _T_2071; // @[AesSbox.scala 40:63]
  wire  _T_2095 = _T_2077 ^ _T_2087; // @[AesSbox.scala 40:63]
  wire  _T_2097 = _T_2089 ^ _T_2083; // @[AesSbox.scala 40:63]
  wire  _T_2099 = _T_2091 ^ _T_2087; // @[AesSbox.scala 40:63]
  wire  _T_2101 = _T_2093 ^ _T_2083; // @[AesSbox.scala 40:63]
  wire  _T_2103 = _T_2095 ^ _T_2025; // @[AesSbox.scala 40:63]
  wire  _T_2105 = _T_2101 ^ _T_2103; // @[AesSbox.scala 40:63]
  wire  _T_2107 = _T_2101 & _T_2097; // @[AesSbox.scala 41:63]
  wire  _T_2109 = _T_2099 ^ _T_2107; // @[AesSbox.scala 40:63]
  wire  _T_2111 = _T_2097 ^ _T_2099; // @[AesSbox.scala 40:63]
  wire  _T_2113 = _T_2103 ^ _T_2107; // @[AesSbox.scala 40:63]
  wire  _T_2115 = _T_2113 & _T_2111; // @[AesSbox.scala 41:63]
  wire  _T_2117 = _T_2109 & _T_2105; // @[AesSbox.scala 41:63]
  wire  _T_2119 = _T_2097 & _T_2103; // @[AesSbox.scala 41:63]
  wire  _T_2121 = _T_2111 & _T_2119; // @[AesSbox.scala 41:63]
  wire  _T_2123 = _T_2111 ^ _T_2107; // @[AesSbox.scala 40:63]
  wire  _T_2125 = _T_2099 & _T_2101; // @[AesSbox.scala 41:63]
  wire  _T_2127 = _T_2105 & _T_2125; // @[AesSbox.scala 41:63]
  wire  _T_2129 = _T_2105 ^ _T_2107; // @[AesSbox.scala 40:63]
  wire  _T_2131 = _T_2099 ^ _T_2115; // @[AesSbox.scala 40:63]
  wire  _T_2133 = _T_2121 ^ _T_2123; // @[AesSbox.scala 40:63]
  wire  _T_2135 = _T_2103 ^ _T_2117; // @[AesSbox.scala 40:63]
  wire  _T_2137 = _T_2127 ^ _T_2129; // @[AesSbox.scala 40:63]
  wire  _T_2139 = _T_2133 ^ _T_2137; // @[AesSbox.scala 40:63]
  wire  _T_2141 = _T_2131 ^ _T_2135; // @[AesSbox.scala 40:63]
  wire  _T_2143 = _T_2131 ^ _T_2133; // @[AesSbox.scala 40:63]
  wire  _T_2145 = _T_2135 ^ _T_2137; // @[AesSbox.scala 40:63]
  wire  _T_2147 = _T_2141 ^ _T_2139; // @[AesSbox.scala 40:63]
  wire  _T_2149 = _T_2145 & _T_2047; // @[AesSbox.scala 41:63]
  wire  _T_2151 = _T_2137 & _T_2011; // @[AesSbox.scala 41:63]
  wire  _T_2153 = _T_2135 & _T_2045; // @[AesSbox.scala 41:63]
  wire  _T_2155 = _T_2143 & _T_2049; // @[AesSbox.scala 41:63]
  wire  _T_2157 = _T_2133 & _T_2016; // @[AesSbox.scala 41:63]
  wire  _T_2159 = _T_2131 & _T_2030; // @[AesSbox.scala 41:63]
  wire  _T_2161 = _T_2141 & _T_2053; // @[AesSbox.scala 41:63]
  wire  _T_2163 = _T_2147 & _T_2051; // @[AesSbox.scala 41:63]
  wire  _T_2165 = _T_2139 & _T_2018; // @[AesSbox.scala 41:63]
  wire  _T_2167 = _T_2145 & _T_2020; // @[AesSbox.scala 41:63]
  wire  _T_2169 = _T_2137 & _T_1995; // @[AesSbox.scala 41:63]
  wire  _T_2171 = _T_2135 & _T_2013; // @[AesSbox.scala 41:63]
  wire  _T_2173 = _T_2143 & _T_2022; // @[AesSbox.scala 41:63]
  wire  _T_2175 = _T_2133 & _T_1998; // @[AesSbox.scala 41:63]
  wire  _T_2177 = _T_2131 & _T_2032; // @[AesSbox.scala 41:63]
  wire  _T_2179 = _T_2141 & _T_2003; // @[AesSbox.scala 41:63]
  wire  _T_2181 = _T_2147 & _T_2034; // @[AesSbox.scala 41:63]
  wire  _T_2183 = _T_2139 & _T_2001; // @[AesSbox.scala 41:63]
  wire  _T_2185 = _T_2161 ^ _T_2179; // @[AesSbox.scala 40:63]
  wire  _T_2187 = _T_2173 ^ _T_2175; // @[AesSbox.scala 40:63]
  wire  _T_2189 = _T_2165 ^ _T_2181; // @[AesSbox.scala 40:63]
  wire  _T_2191 = _T_2151 ^ _T_2157; // @[AesSbox.scala 40:63]
  wire  _T_2193 = _T_2153 ^ _T_2169; // @[AesSbox.scala 40:63]
  wire  _T_2195 = _T_2149 ^ _T_2159; // @[AesSbox.scala 40:63]
  wire  _T_2197 = _T_2155 ^ _T_2177; // @[AesSbox.scala 40:63]
  wire  _T_2199 = _T_2185 ^ _T_2187; // @[AesSbox.scala 40:63]
  wire  _T_2201 = _T_2157 ^ _T_2163; // @[AesSbox.scala 40:63]
  wire  _T_2203 = _T_2167 ^ _T_2183; // @[AesSbox.scala 40:63]
  wire  _T_2205 = _T_2171 ^ _T_2193; // @[AesSbox.scala 40:63]
  wire  _T_2207 = _T_2185 ^ _T_2191; // @[AesSbox.scala 40:63]
  wire  _T_2209 = _T_2149 ^ _T_2153; // @[AesSbox.scala 40:63]
  wire  _T_2211 = _T_2155 ^ _T_2159; // @[AesSbox.scala 40:63]
  wire  _T_2213 = _T_2155 ^ _T_2181; // @[AesSbox.scala 40:63]
  wire  _T_2215 = _T_2165 ^ _T_2175; // @[AesSbox.scala 40:63]
  wire  _T_2217 = _T_2171 ^ _T_2179; // @[AesSbox.scala 40:63]
  wire  _T_2219 = _T_2173 ^ _T_2189; // @[AesSbox.scala 40:63]
  wire  _T_2221 = _T_2183 ^ _T_2195; // @[AesSbox.scala 40:63]
  wire  _T_2223 = _T_2189 ^ _T_2191; // @[AesSbox.scala 40:63]
  wire  _T_2225 = _T_2193 ^ _T_2197; // @[AesSbox.scala 40:63]
  wire  _T_2227 = _T_2189 ^ _T_2199; // @[AesSbox.scala 40:63]
  wire  _T_2229 = _T_2199 ^ _T_2201; // @[AesSbox.scala 40:63]
  wire  _T_2231 = _T_2195 ^ _T_2199; // @[AesSbox.scala 40:63]
  wire  _T_2233 = _T_2197 ^ _T_2205; // @[AesSbox.scala 40:63]
  wire  _T_2235 = _T_2203 ^ _T_2207; // @[AesSbox.scala 40:63]
  wire  _T_2237 = _T_2205 ^ _T_2221; // @[AesSbox.scala 40:63]
  wire  _T_2239 = _T_2207 ^ _T_2233; // @[AesSbox.scala 40:63]
  wire  _T_2241 = _T_2215 ^ _T_2225; // @[AesSbox.scala 40:63]
  wire  _T_2242 = _T_2211 ^ _T_2227; // @[AesSbox.scala 40:63]
  wire  _T_2243 = _T_2235 ^ _T_2241; // @[AesSbox.scala 40:63]
  wire  _T_2244 = _T_2219 ^ _T_2239; // @[AesSbox.scala 40:63]
  wire  _T_2245 = _T_2209 ^ _T_2227; // @[AesSbox.scala 40:63]
  wire  _T_2246 = _T_2229 ^ _T_2237; // @[AesSbox.scala 40:63]
  wire  _T_2247 = _T_2223 ^ _T_2231; // @[AesSbox.scala 40:63]
  wire  _T_2248 = _T_2213 ^ _T_2229; // @[AesSbox.scala 40:63]
  wire  _T_2249 = _T_2203 ^ _T_2217; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_1_3 = {_T_2242,_T_2243,_T_2244,_T_2245,_T_2246,_T_2247,_T_2248,_T_2249}; // @[Cat.scala 29:58]
  wire  _T_2275 = matrix_2_0[7] ^ matrix_2_0[4]; // @[AesSbox.scala 40:63]
  wire  _T_2277 = matrix_2_0[6] ^ matrix_2_0[4]; // @[AesSbox.scala 42:65]
  wire  _T_2278 = ~_T_2277; // @[AesSbox.scala 42:51]
  wire  _T_2280 = matrix_2_0[7] ^ matrix_2_0[6]; // @[AesSbox.scala 42:65]
  wire  _T_2281 = ~_T_2280; // @[AesSbox.scala 42:51]
  wire  _T_2283 = matrix_2_0[4] ^ matrix_2_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_2285 = matrix_2_0[3] ^ matrix_2_0[0]; // @[AesSbox.scala 42:65]
  wire  _T_2286 = ~_T_2285; // @[AesSbox.scala 42:51]
  wire  _T_2288 = matrix_2_0[1] ^ matrix_2_0[0]; // @[AesSbox.scala 40:63]
  wire  _T_2290 = matrix_2_0[6] ^ _T_2275; // @[AesSbox.scala 42:65]
  wire  _T_2291 = ~_T_2290; // @[AesSbox.scala 42:51]
  wire  _T_2293 = _T_2278 ^ _T_2288; // @[AesSbox.scala 40:63]
  wire  _T_2295 = matrix_2_0[0] ^ _T_2283; // @[AesSbox.scala 42:65]
  wire  _T_2296 = ~_T_2295; // @[AesSbox.scala 42:51]
  wire  _T_2298 = _T_2281 ^ _T_2286; // @[AesSbox.scala 40:63]
  wire  _T_2300 = _T_2281 ^ _T_2288; // @[AesSbox.scala 40:63]
  wire  _T_2302 = _T_2283 ^ _T_2288; // @[AesSbox.scala 40:63]
  wire  _T_2304 = matrix_2_0[5] ^ _T_2283; // @[AesSbox.scala 42:65]
  wire  _T_2305 = ~_T_2304; // @[AesSbox.scala 42:51]
  wire  _T_2307 = matrix_2_0[6] ^ matrix_2_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_2309 = matrix_2_0[5] ^ _T_2293; // @[AesSbox.scala 42:65]
  wire  _T_2310 = ~_T_2309; // @[AesSbox.scala 42:51]
  wire  _T_2312 = _T_2286 ^ _T_2307; // @[AesSbox.scala 40:63]
  wire  _T_2314 = matrix_2_0[3] ^ _T_2291; // @[AesSbox.scala 40:63]
  wire  _T_2316 = matrix_2_0[5] ^ matrix_2_0[2]; // @[AesSbox.scala 42:65]
  wire  _T_2317 = ~_T_2316; // @[AesSbox.scala 42:51]
  wire  _T_2319 = matrix_2_0[2] ^ matrix_2_0[1]; // @[AesSbox.scala 42:65]
  wire  _T_2320 = ~_T_2319; // @[AesSbox.scala 42:51]
  wire  _T_2322 = matrix_2_0[5] ^ matrix_2_0[3]; // @[AesSbox.scala 42:65]
  wire  _T_2323 = ~_T_2322; // @[AesSbox.scala 42:51]
  wire  _T_2325 = matrix_2_0[7] ^ _T_2317; // @[AesSbox.scala 40:63]
  wire  _T_2327 = _T_2278 ^ _T_2317; // @[AesSbox.scala 40:63]
  wire  _T_2329 = _T_2307 ^ _T_2323; // @[AesSbox.scala 40:63]
  wire  _T_2331 = _T_2283 ^ _T_2320; // @[AesSbox.scala 40:63]
  wire  _T_2333 = _T_2298 ^ _T_2331; // @[AesSbox.scala 40:63]
  wire  _T_2335 = _T_2298 ^ _T_2320; // @[AesSbox.scala 40:63]
  wire  _T_2337 = _T_2302 ^ _T_2329; // @[AesSbox.scala 40:63]
  wire  _T_2339 = _T_2300 & _T_2327; // @[AesSbox.scala 41:63]
  wire  _T_2341 = _T_2275 & _T_2291; // @[AesSbox.scala 41:63]
  wire  _T_2343 = _T_2335 ^ _T_2339; // @[AesSbox.scala 40:63]
  wire  _T_2345 = _T_2293 & _T_2325; // @[AesSbox.scala 41:63]
  wire  _T_2347 = _T_2345 ^ _T_2339; // @[AesSbox.scala 40:63]
  wire  _T_2349 = _T_2302 & _T_2329; // @[AesSbox.scala 41:63]
  wire  _T_2351 = _T_2278 & _T_2296; // @[AesSbox.scala 41:63]
  wire  _T_2353 = _T_2337 ^ _T_2349; // @[AesSbox.scala 40:63]
  wire  _T_2355 = _T_2312 & _T_2310; // @[AesSbox.scala 41:63]
  wire  _T_2357 = _T_2355 ^ _T_2349; // @[AesSbox.scala 40:63]
  wire  _T_2359 = _T_2283 & _T_2333; // @[AesSbox.scala 41:63]
  wire  _T_2361 = _T_2314 & _T_2331; // @[AesSbox.scala 41:63]
  wire  _T_2363 = _T_2361 ^ _T_2359; // @[AesSbox.scala 40:63]
  wire  _T_2365 = _T_2281 & _T_2298; // @[AesSbox.scala 41:63]
  wire  _T_2367 = _T_2365 ^ _T_2359; // @[AesSbox.scala 40:63]
  wire  _T_2369 = _T_2343 ^ _T_2341; // @[AesSbox.scala 40:63]
  wire  _T_2371 = _T_2347 ^ _T_2286; // @[AesSbox.scala 40:63]
  wire  _T_2373 = _T_2353 ^ _T_2351; // @[AesSbox.scala 40:63]
  wire  _T_2375 = _T_2357 ^ _T_2367; // @[AesSbox.scala 40:63]
  wire  _T_2377 = _T_2369 ^ _T_2363; // @[AesSbox.scala 40:63]
  wire  _T_2379 = _T_2371 ^ _T_2367; // @[AesSbox.scala 40:63]
  wire  _T_2381 = _T_2373 ^ _T_2363; // @[AesSbox.scala 40:63]
  wire  _T_2383 = _T_2375 ^ _T_2305; // @[AesSbox.scala 40:63]
  wire  _T_2385 = _T_2381 ^ _T_2383; // @[AesSbox.scala 40:63]
  wire  _T_2387 = _T_2381 & _T_2377; // @[AesSbox.scala 41:63]
  wire  _T_2389 = _T_2379 ^ _T_2387; // @[AesSbox.scala 40:63]
  wire  _T_2391 = _T_2377 ^ _T_2379; // @[AesSbox.scala 40:63]
  wire  _T_2393 = _T_2383 ^ _T_2387; // @[AesSbox.scala 40:63]
  wire  _T_2395 = _T_2393 & _T_2391; // @[AesSbox.scala 41:63]
  wire  _T_2397 = _T_2389 & _T_2385; // @[AesSbox.scala 41:63]
  wire  _T_2399 = _T_2377 & _T_2383; // @[AesSbox.scala 41:63]
  wire  _T_2401 = _T_2391 & _T_2399; // @[AesSbox.scala 41:63]
  wire  _T_2403 = _T_2391 ^ _T_2387; // @[AesSbox.scala 40:63]
  wire  _T_2405 = _T_2379 & _T_2381; // @[AesSbox.scala 41:63]
  wire  _T_2407 = _T_2385 & _T_2405; // @[AesSbox.scala 41:63]
  wire  _T_2409 = _T_2385 ^ _T_2387; // @[AesSbox.scala 40:63]
  wire  _T_2411 = _T_2379 ^ _T_2395; // @[AesSbox.scala 40:63]
  wire  _T_2413 = _T_2401 ^ _T_2403; // @[AesSbox.scala 40:63]
  wire  _T_2415 = _T_2383 ^ _T_2397; // @[AesSbox.scala 40:63]
  wire  _T_2417 = _T_2407 ^ _T_2409; // @[AesSbox.scala 40:63]
  wire  _T_2419 = _T_2413 ^ _T_2417; // @[AesSbox.scala 40:63]
  wire  _T_2421 = _T_2411 ^ _T_2415; // @[AesSbox.scala 40:63]
  wire  _T_2423 = _T_2411 ^ _T_2413; // @[AesSbox.scala 40:63]
  wire  _T_2425 = _T_2415 ^ _T_2417; // @[AesSbox.scala 40:63]
  wire  _T_2427 = _T_2421 ^ _T_2419; // @[AesSbox.scala 40:63]
  wire  _T_2429 = _T_2425 & _T_2327; // @[AesSbox.scala 41:63]
  wire  _T_2431 = _T_2417 & _T_2291; // @[AesSbox.scala 41:63]
  wire  _T_2433 = _T_2415 & _T_2325; // @[AesSbox.scala 41:63]
  wire  _T_2435 = _T_2423 & _T_2329; // @[AesSbox.scala 41:63]
  wire  _T_2437 = _T_2413 & _T_2296; // @[AesSbox.scala 41:63]
  wire  _T_2439 = _T_2411 & _T_2310; // @[AesSbox.scala 41:63]
  wire  _T_2441 = _T_2421 & _T_2333; // @[AesSbox.scala 41:63]
  wire  _T_2443 = _T_2427 & _T_2331; // @[AesSbox.scala 41:63]
  wire  _T_2445 = _T_2419 & _T_2298; // @[AesSbox.scala 41:63]
  wire  _T_2447 = _T_2425 & _T_2300; // @[AesSbox.scala 41:63]
  wire  _T_2449 = _T_2417 & _T_2275; // @[AesSbox.scala 41:63]
  wire  _T_2451 = _T_2415 & _T_2293; // @[AesSbox.scala 41:63]
  wire  _T_2453 = _T_2423 & _T_2302; // @[AesSbox.scala 41:63]
  wire  _T_2455 = _T_2413 & _T_2278; // @[AesSbox.scala 41:63]
  wire  _T_2457 = _T_2411 & _T_2312; // @[AesSbox.scala 41:63]
  wire  _T_2459 = _T_2421 & _T_2283; // @[AesSbox.scala 41:63]
  wire  _T_2461 = _T_2427 & _T_2314; // @[AesSbox.scala 41:63]
  wire  _T_2463 = _T_2419 & _T_2281; // @[AesSbox.scala 41:63]
  wire  _T_2465 = _T_2441 ^ _T_2459; // @[AesSbox.scala 40:63]
  wire  _T_2467 = _T_2453 ^ _T_2455; // @[AesSbox.scala 40:63]
  wire  _T_2469 = _T_2445 ^ _T_2461; // @[AesSbox.scala 40:63]
  wire  _T_2471 = _T_2431 ^ _T_2437; // @[AesSbox.scala 40:63]
  wire  _T_2473 = _T_2433 ^ _T_2449; // @[AesSbox.scala 40:63]
  wire  _T_2475 = _T_2429 ^ _T_2439; // @[AesSbox.scala 40:63]
  wire  _T_2477 = _T_2435 ^ _T_2457; // @[AesSbox.scala 40:63]
  wire  _T_2479 = _T_2465 ^ _T_2467; // @[AesSbox.scala 40:63]
  wire  _T_2481 = _T_2437 ^ _T_2443; // @[AesSbox.scala 40:63]
  wire  _T_2483 = _T_2447 ^ _T_2463; // @[AesSbox.scala 40:63]
  wire  _T_2485 = _T_2451 ^ _T_2473; // @[AesSbox.scala 40:63]
  wire  _T_2487 = _T_2465 ^ _T_2471; // @[AesSbox.scala 40:63]
  wire  _T_2489 = _T_2429 ^ _T_2433; // @[AesSbox.scala 40:63]
  wire  _T_2491 = _T_2435 ^ _T_2439; // @[AesSbox.scala 40:63]
  wire  _T_2493 = _T_2435 ^ _T_2461; // @[AesSbox.scala 40:63]
  wire  _T_2495 = _T_2445 ^ _T_2455; // @[AesSbox.scala 40:63]
  wire  _T_2497 = _T_2451 ^ _T_2459; // @[AesSbox.scala 40:63]
  wire  _T_2499 = _T_2453 ^ _T_2469; // @[AesSbox.scala 40:63]
  wire  _T_2501 = _T_2463 ^ _T_2475; // @[AesSbox.scala 40:63]
  wire  _T_2503 = _T_2469 ^ _T_2471; // @[AesSbox.scala 40:63]
  wire  _T_2505 = _T_2473 ^ _T_2477; // @[AesSbox.scala 40:63]
  wire  _T_2507 = _T_2469 ^ _T_2479; // @[AesSbox.scala 40:63]
  wire  _T_2509 = _T_2479 ^ _T_2481; // @[AesSbox.scala 40:63]
  wire  _T_2511 = _T_2475 ^ _T_2479; // @[AesSbox.scala 40:63]
  wire  _T_2513 = _T_2477 ^ _T_2485; // @[AesSbox.scala 40:63]
  wire  _T_2515 = _T_2483 ^ _T_2487; // @[AesSbox.scala 40:63]
  wire  _T_2517 = _T_2485 ^ _T_2501; // @[AesSbox.scala 40:63]
  wire  _T_2519 = _T_2487 ^ _T_2513; // @[AesSbox.scala 40:63]
  wire  _T_2521 = _T_2495 ^ _T_2505; // @[AesSbox.scala 40:63]
  wire  _T_2522 = _T_2491 ^ _T_2507; // @[AesSbox.scala 40:63]
  wire  _T_2523 = _T_2515 ^ _T_2521; // @[AesSbox.scala 40:63]
  wire  _T_2524 = _T_2499 ^ _T_2519; // @[AesSbox.scala 40:63]
  wire  _T_2525 = _T_2489 ^ _T_2507; // @[AesSbox.scala 40:63]
  wire  _T_2526 = _T_2509 ^ _T_2517; // @[AesSbox.scala 40:63]
  wire  _T_2527 = _T_2503 ^ _T_2511; // @[AesSbox.scala 40:63]
  wire  _T_2528 = _T_2493 ^ _T_2509; // @[AesSbox.scala 40:63]
  wire  _T_2529 = _T_2483 ^ _T_2497; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_2_0 = {_T_2522,_T_2523,_T_2524,_T_2525,_T_2526,_T_2527,_T_2528,_T_2529}; // @[Cat.scala 29:58]
  wire  _T_2554 = matrix_1_1[7] ^ matrix_1_1[4]; // @[AesSbox.scala 40:63]
  wire  _T_2556 = matrix_1_1[6] ^ matrix_1_1[4]; // @[AesSbox.scala 42:65]
  wire  _T_2557 = ~_T_2556; // @[AesSbox.scala 42:51]
  wire  _T_2559 = matrix_1_1[7] ^ matrix_1_1[6]; // @[AesSbox.scala 42:65]
  wire  _T_2560 = ~_T_2559; // @[AesSbox.scala 42:51]
  wire  _T_2562 = matrix_1_1[4] ^ matrix_1_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_2564 = matrix_1_1[3] ^ matrix_1_1[0]; // @[AesSbox.scala 42:65]
  wire  _T_2565 = ~_T_2564; // @[AesSbox.scala 42:51]
  wire  _T_2567 = matrix_1_1[1] ^ matrix_1_1[0]; // @[AesSbox.scala 40:63]
  wire  _T_2569 = matrix_1_1[6] ^ _T_2554; // @[AesSbox.scala 42:65]
  wire  _T_2570 = ~_T_2569; // @[AesSbox.scala 42:51]
  wire  _T_2572 = _T_2557 ^ _T_2567; // @[AesSbox.scala 40:63]
  wire  _T_2574 = matrix_1_1[0] ^ _T_2562; // @[AesSbox.scala 42:65]
  wire  _T_2575 = ~_T_2574; // @[AesSbox.scala 42:51]
  wire  _T_2577 = _T_2560 ^ _T_2565; // @[AesSbox.scala 40:63]
  wire  _T_2579 = _T_2560 ^ _T_2567; // @[AesSbox.scala 40:63]
  wire  _T_2581 = _T_2562 ^ _T_2567; // @[AesSbox.scala 40:63]
  wire  _T_2583 = matrix_1_1[5] ^ _T_2562; // @[AesSbox.scala 42:65]
  wire  _T_2584 = ~_T_2583; // @[AesSbox.scala 42:51]
  wire  _T_2586 = matrix_1_1[6] ^ matrix_1_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_2588 = matrix_1_1[5] ^ _T_2572; // @[AesSbox.scala 42:65]
  wire  _T_2589 = ~_T_2588; // @[AesSbox.scala 42:51]
  wire  _T_2591 = _T_2565 ^ _T_2586; // @[AesSbox.scala 40:63]
  wire  _T_2593 = matrix_1_1[3] ^ _T_2570; // @[AesSbox.scala 40:63]
  wire  _T_2595 = matrix_1_1[5] ^ matrix_1_1[2]; // @[AesSbox.scala 42:65]
  wire  _T_2596 = ~_T_2595; // @[AesSbox.scala 42:51]
  wire  _T_2598 = matrix_1_1[2] ^ matrix_1_1[1]; // @[AesSbox.scala 42:65]
  wire  _T_2599 = ~_T_2598; // @[AesSbox.scala 42:51]
  wire  _T_2601 = matrix_1_1[5] ^ matrix_1_1[3]; // @[AesSbox.scala 42:65]
  wire  _T_2602 = ~_T_2601; // @[AesSbox.scala 42:51]
  wire  _T_2604 = matrix_1_1[7] ^ _T_2596; // @[AesSbox.scala 40:63]
  wire  _T_2606 = _T_2557 ^ _T_2596; // @[AesSbox.scala 40:63]
  wire  _T_2608 = _T_2586 ^ _T_2602; // @[AesSbox.scala 40:63]
  wire  _T_2610 = _T_2562 ^ _T_2599; // @[AesSbox.scala 40:63]
  wire  _T_2612 = _T_2577 ^ _T_2610; // @[AesSbox.scala 40:63]
  wire  _T_2614 = _T_2577 ^ _T_2599; // @[AesSbox.scala 40:63]
  wire  _T_2616 = _T_2581 ^ _T_2608; // @[AesSbox.scala 40:63]
  wire  _T_2618 = _T_2579 & _T_2606; // @[AesSbox.scala 41:63]
  wire  _T_2620 = _T_2554 & _T_2570; // @[AesSbox.scala 41:63]
  wire  _T_2622 = _T_2614 ^ _T_2618; // @[AesSbox.scala 40:63]
  wire  _T_2624 = _T_2572 & _T_2604; // @[AesSbox.scala 41:63]
  wire  _T_2626 = _T_2624 ^ _T_2618; // @[AesSbox.scala 40:63]
  wire  _T_2628 = _T_2581 & _T_2608; // @[AesSbox.scala 41:63]
  wire  _T_2630 = _T_2557 & _T_2575; // @[AesSbox.scala 41:63]
  wire  _T_2632 = _T_2616 ^ _T_2628; // @[AesSbox.scala 40:63]
  wire  _T_2634 = _T_2591 & _T_2589; // @[AesSbox.scala 41:63]
  wire  _T_2636 = _T_2634 ^ _T_2628; // @[AesSbox.scala 40:63]
  wire  _T_2638 = _T_2562 & _T_2612; // @[AesSbox.scala 41:63]
  wire  _T_2640 = _T_2593 & _T_2610; // @[AesSbox.scala 41:63]
  wire  _T_2642 = _T_2640 ^ _T_2638; // @[AesSbox.scala 40:63]
  wire  _T_2644 = _T_2560 & _T_2577; // @[AesSbox.scala 41:63]
  wire  _T_2646 = _T_2644 ^ _T_2638; // @[AesSbox.scala 40:63]
  wire  _T_2648 = _T_2622 ^ _T_2620; // @[AesSbox.scala 40:63]
  wire  _T_2650 = _T_2626 ^ _T_2565; // @[AesSbox.scala 40:63]
  wire  _T_2652 = _T_2632 ^ _T_2630; // @[AesSbox.scala 40:63]
  wire  _T_2654 = _T_2636 ^ _T_2646; // @[AesSbox.scala 40:63]
  wire  _T_2656 = _T_2648 ^ _T_2642; // @[AesSbox.scala 40:63]
  wire  _T_2658 = _T_2650 ^ _T_2646; // @[AesSbox.scala 40:63]
  wire  _T_2660 = _T_2652 ^ _T_2642; // @[AesSbox.scala 40:63]
  wire  _T_2662 = _T_2654 ^ _T_2584; // @[AesSbox.scala 40:63]
  wire  _T_2664 = _T_2660 ^ _T_2662; // @[AesSbox.scala 40:63]
  wire  _T_2666 = _T_2660 & _T_2656; // @[AesSbox.scala 41:63]
  wire  _T_2668 = _T_2658 ^ _T_2666; // @[AesSbox.scala 40:63]
  wire  _T_2670 = _T_2656 ^ _T_2658; // @[AesSbox.scala 40:63]
  wire  _T_2672 = _T_2662 ^ _T_2666; // @[AesSbox.scala 40:63]
  wire  _T_2674 = _T_2672 & _T_2670; // @[AesSbox.scala 41:63]
  wire  _T_2676 = _T_2668 & _T_2664; // @[AesSbox.scala 41:63]
  wire  _T_2678 = _T_2656 & _T_2662; // @[AesSbox.scala 41:63]
  wire  _T_2680 = _T_2670 & _T_2678; // @[AesSbox.scala 41:63]
  wire  _T_2682 = _T_2670 ^ _T_2666; // @[AesSbox.scala 40:63]
  wire  _T_2684 = _T_2658 & _T_2660; // @[AesSbox.scala 41:63]
  wire  _T_2686 = _T_2664 & _T_2684; // @[AesSbox.scala 41:63]
  wire  _T_2688 = _T_2664 ^ _T_2666; // @[AesSbox.scala 40:63]
  wire  _T_2690 = _T_2658 ^ _T_2674; // @[AesSbox.scala 40:63]
  wire  _T_2692 = _T_2680 ^ _T_2682; // @[AesSbox.scala 40:63]
  wire  _T_2694 = _T_2662 ^ _T_2676; // @[AesSbox.scala 40:63]
  wire  _T_2696 = _T_2686 ^ _T_2688; // @[AesSbox.scala 40:63]
  wire  _T_2698 = _T_2692 ^ _T_2696; // @[AesSbox.scala 40:63]
  wire  _T_2700 = _T_2690 ^ _T_2694; // @[AesSbox.scala 40:63]
  wire  _T_2702 = _T_2690 ^ _T_2692; // @[AesSbox.scala 40:63]
  wire  _T_2704 = _T_2694 ^ _T_2696; // @[AesSbox.scala 40:63]
  wire  _T_2706 = _T_2700 ^ _T_2698; // @[AesSbox.scala 40:63]
  wire  _T_2708 = _T_2704 & _T_2606; // @[AesSbox.scala 41:63]
  wire  _T_2710 = _T_2696 & _T_2570; // @[AesSbox.scala 41:63]
  wire  _T_2712 = _T_2694 & _T_2604; // @[AesSbox.scala 41:63]
  wire  _T_2714 = _T_2702 & _T_2608; // @[AesSbox.scala 41:63]
  wire  _T_2716 = _T_2692 & _T_2575; // @[AesSbox.scala 41:63]
  wire  _T_2718 = _T_2690 & _T_2589; // @[AesSbox.scala 41:63]
  wire  _T_2720 = _T_2700 & _T_2612; // @[AesSbox.scala 41:63]
  wire  _T_2722 = _T_2706 & _T_2610; // @[AesSbox.scala 41:63]
  wire  _T_2724 = _T_2698 & _T_2577; // @[AesSbox.scala 41:63]
  wire  _T_2726 = _T_2704 & _T_2579; // @[AesSbox.scala 41:63]
  wire  _T_2728 = _T_2696 & _T_2554; // @[AesSbox.scala 41:63]
  wire  _T_2730 = _T_2694 & _T_2572; // @[AesSbox.scala 41:63]
  wire  _T_2732 = _T_2702 & _T_2581; // @[AesSbox.scala 41:63]
  wire  _T_2734 = _T_2692 & _T_2557; // @[AesSbox.scala 41:63]
  wire  _T_2736 = _T_2690 & _T_2591; // @[AesSbox.scala 41:63]
  wire  _T_2738 = _T_2700 & _T_2562; // @[AesSbox.scala 41:63]
  wire  _T_2740 = _T_2706 & _T_2593; // @[AesSbox.scala 41:63]
  wire  _T_2742 = _T_2698 & _T_2560; // @[AesSbox.scala 41:63]
  wire  _T_2744 = _T_2720 ^ _T_2738; // @[AesSbox.scala 40:63]
  wire  _T_2746 = _T_2732 ^ _T_2734; // @[AesSbox.scala 40:63]
  wire  _T_2748 = _T_2724 ^ _T_2740; // @[AesSbox.scala 40:63]
  wire  _T_2750 = _T_2710 ^ _T_2716; // @[AesSbox.scala 40:63]
  wire  _T_2752 = _T_2712 ^ _T_2728; // @[AesSbox.scala 40:63]
  wire  _T_2754 = _T_2708 ^ _T_2718; // @[AesSbox.scala 40:63]
  wire  _T_2756 = _T_2714 ^ _T_2736; // @[AesSbox.scala 40:63]
  wire  _T_2758 = _T_2744 ^ _T_2746; // @[AesSbox.scala 40:63]
  wire  _T_2760 = _T_2716 ^ _T_2722; // @[AesSbox.scala 40:63]
  wire  _T_2762 = _T_2726 ^ _T_2742; // @[AesSbox.scala 40:63]
  wire  _T_2764 = _T_2730 ^ _T_2752; // @[AesSbox.scala 40:63]
  wire  _T_2766 = _T_2744 ^ _T_2750; // @[AesSbox.scala 40:63]
  wire  _T_2768 = _T_2708 ^ _T_2712; // @[AesSbox.scala 40:63]
  wire  _T_2770 = _T_2714 ^ _T_2718; // @[AesSbox.scala 40:63]
  wire  _T_2772 = _T_2714 ^ _T_2740; // @[AesSbox.scala 40:63]
  wire  _T_2774 = _T_2724 ^ _T_2734; // @[AesSbox.scala 40:63]
  wire  _T_2776 = _T_2730 ^ _T_2738; // @[AesSbox.scala 40:63]
  wire  _T_2778 = _T_2732 ^ _T_2748; // @[AesSbox.scala 40:63]
  wire  _T_2780 = _T_2742 ^ _T_2754; // @[AesSbox.scala 40:63]
  wire  _T_2782 = _T_2748 ^ _T_2750; // @[AesSbox.scala 40:63]
  wire  _T_2784 = _T_2752 ^ _T_2756; // @[AesSbox.scala 40:63]
  wire  _T_2786 = _T_2748 ^ _T_2758; // @[AesSbox.scala 40:63]
  wire  _T_2788 = _T_2758 ^ _T_2760; // @[AesSbox.scala 40:63]
  wire  _T_2790 = _T_2754 ^ _T_2758; // @[AesSbox.scala 40:63]
  wire  _T_2792 = _T_2756 ^ _T_2764; // @[AesSbox.scala 40:63]
  wire  _T_2794 = _T_2762 ^ _T_2766; // @[AesSbox.scala 40:63]
  wire  _T_2796 = _T_2764 ^ _T_2780; // @[AesSbox.scala 40:63]
  wire  _T_2798 = _T_2766 ^ _T_2792; // @[AesSbox.scala 40:63]
  wire  _T_2800 = _T_2774 ^ _T_2784; // @[AesSbox.scala 40:63]
  wire  _T_2801 = _T_2770 ^ _T_2786; // @[AesSbox.scala 40:63]
  wire  _T_2802 = _T_2794 ^ _T_2800; // @[AesSbox.scala 40:63]
  wire  _T_2803 = _T_2778 ^ _T_2798; // @[AesSbox.scala 40:63]
  wire  _T_2804 = _T_2768 ^ _T_2786; // @[AesSbox.scala 40:63]
  wire  _T_2805 = _T_2788 ^ _T_2796; // @[AesSbox.scala 40:63]
  wire  _T_2806 = _T_2782 ^ _T_2790; // @[AesSbox.scala 40:63]
  wire  _T_2807 = _T_2772 ^ _T_2788; // @[AesSbox.scala 40:63]
  wire  _T_2808 = _T_2762 ^ _T_2776; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_2_1 = {_T_2801,_T_2802,_T_2803,_T_2804,_T_2805,_T_2806,_T_2807,_T_2808}; // @[Cat.scala 29:58]
  wire  _T_2833 = matrix_0_2[7] ^ matrix_0_2[4]; // @[AesSbox.scala 40:63]
  wire  _T_2835 = matrix_0_2[6] ^ matrix_0_2[4]; // @[AesSbox.scala 42:65]
  wire  _T_2836 = ~_T_2835; // @[AesSbox.scala 42:51]
  wire  _T_2838 = matrix_0_2[7] ^ matrix_0_2[6]; // @[AesSbox.scala 42:65]
  wire  _T_2839 = ~_T_2838; // @[AesSbox.scala 42:51]
  wire  _T_2841 = matrix_0_2[4] ^ matrix_0_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_2843 = matrix_0_2[3] ^ matrix_0_2[0]; // @[AesSbox.scala 42:65]
  wire  _T_2844 = ~_T_2843; // @[AesSbox.scala 42:51]
  wire  _T_2846 = matrix_0_2[1] ^ matrix_0_2[0]; // @[AesSbox.scala 40:63]
  wire  _T_2848 = matrix_0_2[6] ^ _T_2833; // @[AesSbox.scala 42:65]
  wire  _T_2849 = ~_T_2848; // @[AesSbox.scala 42:51]
  wire  _T_2851 = _T_2836 ^ _T_2846; // @[AesSbox.scala 40:63]
  wire  _T_2853 = matrix_0_2[0] ^ _T_2841; // @[AesSbox.scala 42:65]
  wire  _T_2854 = ~_T_2853; // @[AesSbox.scala 42:51]
  wire  _T_2856 = _T_2839 ^ _T_2844; // @[AesSbox.scala 40:63]
  wire  _T_2858 = _T_2839 ^ _T_2846; // @[AesSbox.scala 40:63]
  wire  _T_2860 = _T_2841 ^ _T_2846; // @[AesSbox.scala 40:63]
  wire  _T_2862 = matrix_0_2[5] ^ _T_2841; // @[AesSbox.scala 42:65]
  wire  _T_2863 = ~_T_2862; // @[AesSbox.scala 42:51]
  wire  _T_2865 = matrix_0_2[6] ^ matrix_0_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_2867 = matrix_0_2[5] ^ _T_2851; // @[AesSbox.scala 42:65]
  wire  _T_2868 = ~_T_2867; // @[AesSbox.scala 42:51]
  wire  _T_2870 = _T_2844 ^ _T_2865; // @[AesSbox.scala 40:63]
  wire  _T_2872 = matrix_0_2[3] ^ _T_2849; // @[AesSbox.scala 40:63]
  wire  _T_2874 = matrix_0_2[5] ^ matrix_0_2[2]; // @[AesSbox.scala 42:65]
  wire  _T_2875 = ~_T_2874; // @[AesSbox.scala 42:51]
  wire  _T_2877 = matrix_0_2[2] ^ matrix_0_2[1]; // @[AesSbox.scala 42:65]
  wire  _T_2878 = ~_T_2877; // @[AesSbox.scala 42:51]
  wire  _T_2880 = matrix_0_2[5] ^ matrix_0_2[3]; // @[AesSbox.scala 42:65]
  wire  _T_2881 = ~_T_2880; // @[AesSbox.scala 42:51]
  wire  _T_2883 = matrix_0_2[7] ^ _T_2875; // @[AesSbox.scala 40:63]
  wire  _T_2885 = _T_2836 ^ _T_2875; // @[AesSbox.scala 40:63]
  wire  _T_2887 = _T_2865 ^ _T_2881; // @[AesSbox.scala 40:63]
  wire  _T_2889 = _T_2841 ^ _T_2878; // @[AesSbox.scala 40:63]
  wire  _T_2891 = _T_2856 ^ _T_2889; // @[AesSbox.scala 40:63]
  wire  _T_2893 = _T_2856 ^ _T_2878; // @[AesSbox.scala 40:63]
  wire  _T_2895 = _T_2860 ^ _T_2887; // @[AesSbox.scala 40:63]
  wire  _T_2897 = _T_2858 & _T_2885; // @[AesSbox.scala 41:63]
  wire  _T_2899 = _T_2833 & _T_2849; // @[AesSbox.scala 41:63]
  wire  _T_2901 = _T_2893 ^ _T_2897; // @[AesSbox.scala 40:63]
  wire  _T_2903 = _T_2851 & _T_2883; // @[AesSbox.scala 41:63]
  wire  _T_2905 = _T_2903 ^ _T_2897; // @[AesSbox.scala 40:63]
  wire  _T_2907 = _T_2860 & _T_2887; // @[AesSbox.scala 41:63]
  wire  _T_2909 = _T_2836 & _T_2854; // @[AesSbox.scala 41:63]
  wire  _T_2911 = _T_2895 ^ _T_2907; // @[AesSbox.scala 40:63]
  wire  _T_2913 = _T_2870 & _T_2868; // @[AesSbox.scala 41:63]
  wire  _T_2915 = _T_2913 ^ _T_2907; // @[AesSbox.scala 40:63]
  wire  _T_2917 = _T_2841 & _T_2891; // @[AesSbox.scala 41:63]
  wire  _T_2919 = _T_2872 & _T_2889; // @[AesSbox.scala 41:63]
  wire  _T_2921 = _T_2919 ^ _T_2917; // @[AesSbox.scala 40:63]
  wire  _T_2923 = _T_2839 & _T_2856; // @[AesSbox.scala 41:63]
  wire  _T_2925 = _T_2923 ^ _T_2917; // @[AesSbox.scala 40:63]
  wire  _T_2927 = _T_2901 ^ _T_2899; // @[AesSbox.scala 40:63]
  wire  _T_2929 = _T_2905 ^ _T_2844; // @[AesSbox.scala 40:63]
  wire  _T_2931 = _T_2911 ^ _T_2909; // @[AesSbox.scala 40:63]
  wire  _T_2933 = _T_2915 ^ _T_2925; // @[AesSbox.scala 40:63]
  wire  _T_2935 = _T_2927 ^ _T_2921; // @[AesSbox.scala 40:63]
  wire  _T_2937 = _T_2929 ^ _T_2925; // @[AesSbox.scala 40:63]
  wire  _T_2939 = _T_2931 ^ _T_2921; // @[AesSbox.scala 40:63]
  wire  _T_2941 = _T_2933 ^ _T_2863; // @[AesSbox.scala 40:63]
  wire  _T_2943 = _T_2939 ^ _T_2941; // @[AesSbox.scala 40:63]
  wire  _T_2945 = _T_2939 & _T_2935; // @[AesSbox.scala 41:63]
  wire  _T_2947 = _T_2937 ^ _T_2945; // @[AesSbox.scala 40:63]
  wire  _T_2949 = _T_2935 ^ _T_2937; // @[AesSbox.scala 40:63]
  wire  _T_2951 = _T_2941 ^ _T_2945; // @[AesSbox.scala 40:63]
  wire  _T_2953 = _T_2951 & _T_2949; // @[AesSbox.scala 41:63]
  wire  _T_2955 = _T_2947 & _T_2943; // @[AesSbox.scala 41:63]
  wire  _T_2957 = _T_2935 & _T_2941; // @[AesSbox.scala 41:63]
  wire  _T_2959 = _T_2949 & _T_2957; // @[AesSbox.scala 41:63]
  wire  _T_2961 = _T_2949 ^ _T_2945; // @[AesSbox.scala 40:63]
  wire  _T_2963 = _T_2937 & _T_2939; // @[AesSbox.scala 41:63]
  wire  _T_2965 = _T_2943 & _T_2963; // @[AesSbox.scala 41:63]
  wire  _T_2967 = _T_2943 ^ _T_2945; // @[AesSbox.scala 40:63]
  wire  _T_2969 = _T_2937 ^ _T_2953; // @[AesSbox.scala 40:63]
  wire  _T_2971 = _T_2959 ^ _T_2961; // @[AesSbox.scala 40:63]
  wire  _T_2973 = _T_2941 ^ _T_2955; // @[AesSbox.scala 40:63]
  wire  _T_2975 = _T_2965 ^ _T_2967; // @[AesSbox.scala 40:63]
  wire  _T_2977 = _T_2971 ^ _T_2975; // @[AesSbox.scala 40:63]
  wire  _T_2979 = _T_2969 ^ _T_2973; // @[AesSbox.scala 40:63]
  wire  _T_2981 = _T_2969 ^ _T_2971; // @[AesSbox.scala 40:63]
  wire  _T_2983 = _T_2973 ^ _T_2975; // @[AesSbox.scala 40:63]
  wire  _T_2985 = _T_2979 ^ _T_2977; // @[AesSbox.scala 40:63]
  wire  _T_2987 = _T_2983 & _T_2885; // @[AesSbox.scala 41:63]
  wire  _T_2989 = _T_2975 & _T_2849; // @[AesSbox.scala 41:63]
  wire  _T_2991 = _T_2973 & _T_2883; // @[AesSbox.scala 41:63]
  wire  _T_2993 = _T_2981 & _T_2887; // @[AesSbox.scala 41:63]
  wire  _T_2995 = _T_2971 & _T_2854; // @[AesSbox.scala 41:63]
  wire  _T_2997 = _T_2969 & _T_2868; // @[AesSbox.scala 41:63]
  wire  _T_2999 = _T_2979 & _T_2891; // @[AesSbox.scala 41:63]
  wire  _T_3001 = _T_2985 & _T_2889; // @[AesSbox.scala 41:63]
  wire  _T_3003 = _T_2977 & _T_2856; // @[AesSbox.scala 41:63]
  wire  _T_3005 = _T_2983 & _T_2858; // @[AesSbox.scala 41:63]
  wire  _T_3007 = _T_2975 & _T_2833; // @[AesSbox.scala 41:63]
  wire  _T_3009 = _T_2973 & _T_2851; // @[AesSbox.scala 41:63]
  wire  _T_3011 = _T_2981 & _T_2860; // @[AesSbox.scala 41:63]
  wire  _T_3013 = _T_2971 & _T_2836; // @[AesSbox.scala 41:63]
  wire  _T_3015 = _T_2969 & _T_2870; // @[AesSbox.scala 41:63]
  wire  _T_3017 = _T_2979 & _T_2841; // @[AesSbox.scala 41:63]
  wire  _T_3019 = _T_2985 & _T_2872; // @[AesSbox.scala 41:63]
  wire  _T_3021 = _T_2977 & _T_2839; // @[AesSbox.scala 41:63]
  wire  _T_3023 = _T_2999 ^ _T_3017; // @[AesSbox.scala 40:63]
  wire  _T_3025 = _T_3011 ^ _T_3013; // @[AesSbox.scala 40:63]
  wire  _T_3027 = _T_3003 ^ _T_3019; // @[AesSbox.scala 40:63]
  wire  _T_3029 = _T_2989 ^ _T_2995; // @[AesSbox.scala 40:63]
  wire  _T_3031 = _T_2991 ^ _T_3007; // @[AesSbox.scala 40:63]
  wire  _T_3033 = _T_2987 ^ _T_2997; // @[AesSbox.scala 40:63]
  wire  _T_3035 = _T_2993 ^ _T_3015; // @[AesSbox.scala 40:63]
  wire  _T_3037 = _T_3023 ^ _T_3025; // @[AesSbox.scala 40:63]
  wire  _T_3039 = _T_2995 ^ _T_3001; // @[AesSbox.scala 40:63]
  wire  _T_3041 = _T_3005 ^ _T_3021; // @[AesSbox.scala 40:63]
  wire  _T_3043 = _T_3009 ^ _T_3031; // @[AesSbox.scala 40:63]
  wire  _T_3045 = _T_3023 ^ _T_3029; // @[AesSbox.scala 40:63]
  wire  _T_3047 = _T_2987 ^ _T_2991; // @[AesSbox.scala 40:63]
  wire  _T_3049 = _T_2993 ^ _T_2997; // @[AesSbox.scala 40:63]
  wire  _T_3051 = _T_2993 ^ _T_3019; // @[AesSbox.scala 40:63]
  wire  _T_3053 = _T_3003 ^ _T_3013; // @[AesSbox.scala 40:63]
  wire  _T_3055 = _T_3009 ^ _T_3017; // @[AesSbox.scala 40:63]
  wire  _T_3057 = _T_3011 ^ _T_3027; // @[AesSbox.scala 40:63]
  wire  _T_3059 = _T_3021 ^ _T_3033; // @[AesSbox.scala 40:63]
  wire  _T_3061 = _T_3027 ^ _T_3029; // @[AesSbox.scala 40:63]
  wire  _T_3063 = _T_3031 ^ _T_3035; // @[AesSbox.scala 40:63]
  wire  _T_3065 = _T_3027 ^ _T_3037; // @[AesSbox.scala 40:63]
  wire  _T_3067 = _T_3037 ^ _T_3039; // @[AesSbox.scala 40:63]
  wire  _T_3069 = _T_3033 ^ _T_3037; // @[AesSbox.scala 40:63]
  wire  _T_3071 = _T_3035 ^ _T_3043; // @[AesSbox.scala 40:63]
  wire  _T_3073 = _T_3041 ^ _T_3045; // @[AesSbox.scala 40:63]
  wire  _T_3075 = _T_3043 ^ _T_3059; // @[AesSbox.scala 40:63]
  wire  _T_3077 = _T_3045 ^ _T_3071; // @[AesSbox.scala 40:63]
  wire  _T_3079 = _T_3053 ^ _T_3063; // @[AesSbox.scala 40:63]
  wire  _T_3080 = _T_3049 ^ _T_3065; // @[AesSbox.scala 40:63]
  wire  _T_3081 = _T_3073 ^ _T_3079; // @[AesSbox.scala 40:63]
  wire  _T_3082 = _T_3057 ^ _T_3077; // @[AesSbox.scala 40:63]
  wire  _T_3083 = _T_3047 ^ _T_3065; // @[AesSbox.scala 40:63]
  wire  _T_3084 = _T_3067 ^ _T_3075; // @[AesSbox.scala 40:63]
  wire  _T_3085 = _T_3061 ^ _T_3069; // @[AesSbox.scala 40:63]
  wire  _T_3086 = _T_3051 ^ _T_3067; // @[AesSbox.scala 40:63]
  wire  _T_3087 = _T_3041 ^ _T_3055; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_2_2 = {_T_3080,_T_3081,_T_3082,_T_3083,_T_3084,_T_3085,_T_3086,_T_3087}; // @[Cat.scala 29:58]
  wire  _T_3112 = matrix_3_3[7] ^ matrix_3_3[4]; // @[AesSbox.scala 40:63]
  wire  _T_3114 = matrix_3_3[6] ^ matrix_3_3[4]; // @[AesSbox.scala 42:65]
  wire  _T_3115 = ~_T_3114; // @[AesSbox.scala 42:51]
  wire  _T_3117 = matrix_3_3[7] ^ matrix_3_3[6]; // @[AesSbox.scala 42:65]
  wire  _T_3118 = ~_T_3117; // @[AesSbox.scala 42:51]
  wire  _T_3120 = matrix_3_3[4] ^ matrix_3_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_3122 = matrix_3_3[3] ^ matrix_3_3[0]; // @[AesSbox.scala 42:65]
  wire  _T_3123 = ~_T_3122; // @[AesSbox.scala 42:51]
  wire  _T_3125 = matrix_3_3[1] ^ matrix_3_3[0]; // @[AesSbox.scala 40:63]
  wire  _T_3127 = matrix_3_3[6] ^ _T_3112; // @[AesSbox.scala 42:65]
  wire  _T_3128 = ~_T_3127; // @[AesSbox.scala 42:51]
  wire  _T_3130 = _T_3115 ^ _T_3125; // @[AesSbox.scala 40:63]
  wire  _T_3132 = matrix_3_3[0] ^ _T_3120; // @[AesSbox.scala 42:65]
  wire  _T_3133 = ~_T_3132; // @[AesSbox.scala 42:51]
  wire  _T_3135 = _T_3118 ^ _T_3123; // @[AesSbox.scala 40:63]
  wire  _T_3137 = _T_3118 ^ _T_3125; // @[AesSbox.scala 40:63]
  wire  _T_3139 = _T_3120 ^ _T_3125; // @[AesSbox.scala 40:63]
  wire  _T_3141 = matrix_3_3[5] ^ _T_3120; // @[AesSbox.scala 42:65]
  wire  _T_3142 = ~_T_3141; // @[AesSbox.scala 42:51]
  wire  _T_3144 = matrix_3_3[6] ^ matrix_3_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_3146 = matrix_3_3[5] ^ _T_3130; // @[AesSbox.scala 42:65]
  wire  _T_3147 = ~_T_3146; // @[AesSbox.scala 42:51]
  wire  _T_3149 = _T_3123 ^ _T_3144; // @[AesSbox.scala 40:63]
  wire  _T_3151 = matrix_3_3[3] ^ _T_3128; // @[AesSbox.scala 40:63]
  wire  _T_3153 = matrix_3_3[5] ^ matrix_3_3[2]; // @[AesSbox.scala 42:65]
  wire  _T_3154 = ~_T_3153; // @[AesSbox.scala 42:51]
  wire  _T_3156 = matrix_3_3[2] ^ matrix_3_3[1]; // @[AesSbox.scala 42:65]
  wire  _T_3157 = ~_T_3156; // @[AesSbox.scala 42:51]
  wire  _T_3159 = matrix_3_3[5] ^ matrix_3_3[3]; // @[AesSbox.scala 42:65]
  wire  _T_3160 = ~_T_3159; // @[AesSbox.scala 42:51]
  wire  _T_3162 = matrix_3_3[7] ^ _T_3154; // @[AesSbox.scala 40:63]
  wire  _T_3164 = _T_3115 ^ _T_3154; // @[AesSbox.scala 40:63]
  wire  _T_3166 = _T_3144 ^ _T_3160; // @[AesSbox.scala 40:63]
  wire  _T_3168 = _T_3120 ^ _T_3157; // @[AesSbox.scala 40:63]
  wire  _T_3170 = _T_3135 ^ _T_3168; // @[AesSbox.scala 40:63]
  wire  _T_3172 = _T_3135 ^ _T_3157; // @[AesSbox.scala 40:63]
  wire  _T_3174 = _T_3139 ^ _T_3166; // @[AesSbox.scala 40:63]
  wire  _T_3176 = _T_3137 & _T_3164; // @[AesSbox.scala 41:63]
  wire  _T_3178 = _T_3112 & _T_3128; // @[AesSbox.scala 41:63]
  wire  _T_3180 = _T_3172 ^ _T_3176; // @[AesSbox.scala 40:63]
  wire  _T_3182 = _T_3130 & _T_3162; // @[AesSbox.scala 41:63]
  wire  _T_3184 = _T_3182 ^ _T_3176; // @[AesSbox.scala 40:63]
  wire  _T_3186 = _T_3139 & _T_3166; // @[AesSbox.scala 41:63]
  wire  _T_3188 = _T_3115 & _T_3133; // @[AesSbox.scala 41:63]
  wire  _T_3190 = _T_3174 ^ _T_3186; // @[AesSbox.scala 40:63]
  wire  _T_3192 = _T_3149 & _T_3147; // @[AesSbox.scala 41:63]
  wire  _T_3194 = _T_3192 ^ _T_3186; // @[AesSbox.scala 40:63]
  wire  _T_3196 = _T_3120 & _T_3170; // @[AesSbox.scala 41:63]
  wire  _T_3198 = _T_3151 & _T_3168; // @[AesSbox.scala 41:63]
  wire  _T_3200 = _T_3198 ^ _T_3196; // @[AesSbox.scala 40:63]
  wire  _T_3202 = _T_3118 & _T_3135; // @[AesSbox.scala 41:63]
  wire  _T_3204 = _T_3202 ^ _T_3196; // @[AesSbox.scala 40:63]
  wire  _T_3206 = _T_3180 ^ _T_3178; // @[AesSbox.scala 40:63]
  wire  _T_3208 = _T_3184 ^ _T_3123; // @[AesSbox.scala 40:63]
  wire  _T_3210 = _T_3190 ^ _T_3188; // @[AesSbox.scala 40:63]
  wire  _T_3212 = _T_3194 ^ _T_3204; // @[AesSbox.scala 40:63]
  wire  _T_3214 = _T_3206 ^ _T_3200; // @[AesSbox.scala 40:63]
  wire  _T_3216 = _T_3208 ^ _T_3204; // @[AesSbox.scala 40:63]
  wire  _T_3218 = _T_3210 ^ _T_3200; // @[AesSbox.scala 40:63]
  wire  _T_3220 = _T_3212 ^ _T_3142; // @[AesSbox.scala 40:63]
  wire  _T_3222 = _T_3218 ^ _T_3220; // @[AesSbox.scala 40:63]
  wire  _T_3224 = _T_3218 & _T_3214; // @[AesSbox.scala 41:63]
  wire  _T_3226 = _T_3216 ^ _T_3224; // @[AesSbox.scala 40:63]
  wire  _T_3228 = _T_3214 ^ _T_3216; // @[AesSbox.scala 40:63]
  wire  _T_3230 = _T_3220 ^ _T_3224; // @[AesSbox.scala 40:63]
  wire  _T_3232 = _T_3230 & _T_3228; // @[AesSbox.scala 41:63]
  wire  _T_3234 = _T_3226 & _T_3222; // @[AesSbox.scala 41:63]
  wire  _T_3236 = _T_3214 & _T_3220; // @[AesSbox.scala 41:63]
  wire  _T_3238 = _T_3228 & _T_3236; // @[AesSbox.scala 41:63]
  wire  _T_3240 = _T_3228 ^ _T_3224; // @[AesSbox.scala 40:63]
  wire  _T_3242 = _T_3216 & _T_3218; // @[AesSbox.scala 41:63]
  wire  _T_3244 = _T_3222 & _T_3242; // @[AesSbox.scala 41:63]
  wire  _T_3246 = _T_3222 ^ _T_3224; // @[AesSbox.scala 40:63]
  wire  _T_3248 = _T_3216 ^ _T_3232; // @[AesSbox.scala 40:63]
  wire  _T_3250 = _T_3238 ^ _T_3240; // @[AesSbox.scala 40:63]
  wire  _T_3252 = _T_3220 ^ _T_3234; // @[AesSbox.scala 40:63]
  wire  _T_3254 = _T_3244 ^ _T_3246; // @[AesSbox.scala 40:63]
  wire  _T_3256 = _T_3250 ^ _T_3254; // @[AesSbox.scala 40:63]
  wire  _T_3258 = _T_3248 ^ _T_3252; // @[AesSbox.scala 40:63]
  wire  _T_3260 = _T_3248 ^ _T_3250; // @[AesSbox.scala 40:63]
  wire  _T_3262 = _T_3252 ^ _T_3254; // @[AesSbox.scala 40:63]
  wire  _T_3264 = _T_3258 ^ _T_3256; // @[AesSbox.scala 40:63]
  wire  _T_3266 = _T_3262 & _T_3164; // @[AesSbox.scala 41:63]
  wire  _T_3268 = _T_3254 & _T_3128; // @[AesSbox.scala 41:63]
  wire  _T_3270 = _T_3252 & _T_3162; // @[AesSbox.scala 41:63]
  wire  _T_3272 = _T_3260 & _T_3166; // @[AesSbox.scala 41:63]
  wire  _T_3274 = _T_3250 & _T_3133; // @[AesSbox.scala 41:63]
  wire  _T_3276 = _T_3248 & _T_3147; // @[AesSbox.scala 41:63]
  wire  _T_3278 = _T_3258 & _T_3170; // @[AesSbox.scala 41:63]
  wire  _T_3280 = _T_3264 & _T_3168; // @[AesSbox.scala 41:63]
  wire  _T_3282 = _T_3256 & _T_3135; // @[AesSbox.scala 41:63]
  wire  _T_3284 = _T_3262 & _T_3137; // @[AesSbox.scala 41:63]
  wire  _T_3286 = _T_3254 & _T_3112; // @[AesSbox.scala 41:63]
  wire  _T_3288 = _T_3252 & _T_3130; // @[AesSbox.scala 41:63]
  wire  _T_3290 = _T_3260 & _T_3139; // @[AesSbox.scala 41:63]
  wire  _T_3292 = _T_3250 & _T_3115; // @[AesSbox.scala 41:63]
  wire  _T_3294 = _T_3248 & _T_3149; // @[AesSbox.scala 41:63]
  wire  _T_3296 = _T_3258 & _T_3120; // @[AesSbox.scala 41:63]
  wire  _T_3298 = _T_3264 & _T_3151; // @[AesSbox.scala 41:63]
  wire  _T_3300 = _T_3256 & _T_3118; // @[AesSbox.scala 41:63]
  wire  _T_3302 = _T_3278 ^ _T_3296; // @[AesSbox.scala 40:63]
  wire  _T_3304 = _T_3290 ^ _T_3292; // @[AesSbox.scala 40:63]
  wire  _T_3306 = _T_3282 ^ _T_3298; // @[AesSbox.scala 40:63]
  wire  _T_3308 = _T_3268 ^ _T_3274; // @[AesSbox.scala 40:63]
  wire  _T_3310 = _T_3270 ^ _T_3286; // @[AesSbox.scala 40:63]
  wire  _T_3312 = _T_3266 ^ _T_3276; // @[AesSbox.scala 40:63]
  wire  _T_3314 = _T_3272 ^ _T_3294; // @[AesSbox.scala 40:63]
  wire  _T_3316 = _T_3302 ^ _T_3304; // @[AesSbox.scala 40:63]
  wire  _T_3318 = _T_3274 ^ _T_3280; // @[AesSbox.scala 40:63]
  wire  _T_3320 = _T_3284 ^ _T_3300; // @[AesSbox.scala 40:63]
  wire  _T_3322 = _T_3288 ^ _T_3310; // @[AesSbox.scala 40:63]
  wire  _T_3324 = _T_3302 ^ _T_3308; // @[AesSbox.scala 40:63]
  wire  _T_3326 = _T_3266 ^ _T_3270; // @[AesSbox.scala 40:63]
  wire  _T_3328 = _T_3272 ^ _T_3276; // @[AesSbox.scala 40:63]
  wire  _T_3330 = _T_3272 ^ _T_3298; // @[AesSbox.scala 40:63]
  wire  _T_3332 = _T_3282 ^ _T_3292; // @[AesSbox.scala 40:63]
  wire  _T_3334 = _T_3288 ^ _T_3296; // @[AesSbox.scala 40:63]
  wire  _T_3336 = _T_3290 ^ _T_3306; // @[AesSbox.scala 40:63]
  wire  _T_3338 = _T_3300 ^ _T_3312; // @[AesSbox.scala 40:63]
  wire  _T_3340 = _T_3306 ^ _T_3308; // @[AesSbox.scala 40:63]
  wire  _T_3342 = _T_3310 ^ _T_3314; // @[AesSbox.scala 40:63]
  wire  _T_3344 = _T_3306 ^ _T_3316; // @[AesSbox.scala 40:63]
  wire  _T_3346 = _T_3316 ^ _T_3318; // @[AesSbox.scala 40:63]
  wire  _T_3348 = _T_3312 ^ _T_3316; // @[AesSbox.scala 40:63]
  wire  _T_3350 = _T_3314 ^ _T_3322; // @[AesSbox.scala 40:63]
  wire  _T_3352 = _T_3320 ^ _T_3324; // @[AesSbox.scala 40:63]
  wire  _T_3354 = _T_3322 ^ _T_3338; // @[AesSbox.scala 40:63]
  wire  _T_3356 = _T_3324 ^ _T_3350; // @[AesSbox.scala 40:63]
  wire  _T_3358 = _T_3332 ^ _T_3342; // @[AesSbox.scala 40:63]
  wire  _T_3359 = _T_3328 ^ _T_3344; // @[AesSbox.scala 40:63]
  wire  _T_3360 = _T_3352 ^ _T_3358; // @[AesSbox.scala 40:63]
  wire  _T_3361 = _T_3336 ^ _T_3356; // @[AesSbox.scala 40:63]
  wire  _T_3362 = _T_3326 ^ _T_3344; // @[AesSbox.scala 40:63]
  wire  _T_3363 = _T_3346 ^ _T_3354; // @[AesSbox.scala 40:63]
  wire  _T_3364 = _T_3340 ^ _T_3348; // @[AesSbox.scala 40:63]
  wire  _T_3365 = _T_3330 ^ _T_3346; // @[AesSbox.scala 40:63]
  wire  _T_3366 = _T_3320 ^ _T_3334; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_2_3 = {_T_3359,_T_3360,_T_3361,_T_3362,_T_3363,_T_3364,_T_3365,_T_3366}; // @[Cat.scala 29:58]
  wire  _T_3392 = matrix_3_0[7] ^ matrix_3_0[4]; // @[AesSbox.scala 40:63]
  wire  _T_3394 = matrix_3_0[6] ^ matrix_3_0[4]; // @[AesSbox.scala 42:65]
  wire  _T_3395 = ~_T_3394; // @[AesSbox.scala 42:51]
  wire  _T_3397 = matrix_3_0[7] ^ matrix_3_0[6]; // @[AesSbox.scala 42:65]
  wire  _T_3398 = ~_T_3397; // @[AesSbox.scala 42:51]
  wire  _T_3400 = matrix_3_0[4] ^ matrix_3_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_3402 = matrix_3_0[3] ^ matrix_3_0[0]; // @[AesSbox.scala 42:65]
  wire  _T_3403 = ~_T_3402; // @[AesSbox.scala 42:51]
  wire  _T_3405 = matrix_3_0[1] ^ matrix_3_0[0]; // @[AesSbox.scala 40:63]
  wire  _T_3407 = matrix_3_0[6] ^ _T_3392; // @[AesSbox.scala 42:65]
  wire  _T_3408 = ~_T_3407; // @[AesSbox.scala 42:51]
  wire  _T_3410 = _T_3395 ^ _T_3405; // @[AesSbox.scala 40:63]
  wire  _T_3412 = matrix_3_0[0] ^ _T_3400; // @[AesSbox.scala 42:65]
  wire  _T_3413 = ~_T_3412; // @[AesSbox.scala 42:51]
  wire  _T_3415 = _T_3398 ^ _T_3403; // @[AesSbox.scala 40:63]
  wire  _T_3417 = _T_3398 ^ _T_3405; // @[AesSbox.scala 40:63]
  wire  _T_3419 = _T_3400 ^ _T_3405; // @[AesSbox.scala 40:63]
  wire  _T_3421 = matrix_3_0[5] ^ _T_3400; // @[AesSbox.scala 42:65]
  wire  _T_3422 = ~_T_3421; // @[AesSbox.scala 42:51]
  wire  _T_3424 = matrix_3_0[6] ^ matrix_3_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_3426 = matrix_3_0[5] ^ _T_3410; // @[AesSbox.scala 42:65]
  wire  _T_3427 = ~_T_3426; // @[AesSbox.scala 42:51]
  wire  _T_3429 = _T_3403 ^ _T_3424; // @[AesSbox.scala 40:63]
  wire  _T_3431 = matrix_3_0[3] ^ _T_3408; // @[AesSbox.scala 40:63]
  wire  _T_3433 = matrix_3_0[5] ^ matrix_3_0[2]; // @[AesSbox.scala 42:65]
  wire  _T_3434 = ~_T_3433; // @[AesSbox.scala 42:51]
  wire  _T_3436 = matrix_3_0[2] ^ matrix_3_0[1]; // @[AesSbox.scala 42:65]
  wire  _T_3437 = ~_T_3436; // @[AesSbox.scala 42:51]
  wire  _T_3439 = matrix_3_0[5] ^ matrix_3_0[3]; // @[AesSbox.scala 42:65]
  wire  _T_3440 = ~_T_3439; // @[AesSbox.scala 42:51]
  wire  _T_3442 = matrix_3_0[7] ^ _T_3434; // @[AesSbox.scala 40:63]
  wire  _T_3444 = _T_3395 ^ _T_3434; // @[AesSbox.scala 40:63]
  wire  _T_3446 = _T_3424 ^ _T_3440; // @[AesSbox.scala 40:63]
  wire  _T_3448 = _T_3400 ^ _T_3437; // @[AesSbox.scala 40:63]
  wire  _T_3450 = _T_3415 ^ _T_3448; // @[AesSbox.scala 40:63]
  wire  _T_3452 = _T_3415 ^ _T_3437; // @[AesSbox.scala 40:63]
  wire  _T_3454 = _T_3419 ^ _T_3446; // @[AesSbox.scala 40:63]
  wire  _T_3456 = _T_3417 & _T_3444; // @[AesSbox.scala 41:63]
  wire  _T_3458 = _T_3392 & _T_3408; // @[AesSbox.scala 41:63]
  wire  _T_3460 = _T_3452 ^ _T_3456; // @[AesSbox.scala 40:63]
  wire  _T_3462 = _T_3410 & _T_3442; // @[AesSbox.scala 41:63]
  wire  _T_3464 = _T_3462 ^ _T_3456; // @[AesSbox.scala 40:63]
  wire  _T_3466 = _T_3419 & _T_3446; // @[AesSbox.scala 41:63]
  wire  _T_3468 = _T_3395 & _T_3413; // @[AesSbox.scala 41:63]
  wire  _T_3470 = _T_3454 ^ _T_3466; // @[AesSbox.scala 40:63]
  wire  _T_3472 = _T_3429 & _T_3427; // @[AesSbox.scala 41:63]
  wire  _T_3474 = _T_3472 ^ _T_3466; // @[AesSbox.scala 40:63]
  wire  _T_3476 = _T_3400 & _T_3450; // @[AesSbox.scala 41:63]
  wire  _T_3478 = _T_3431 & _T_3448; // @[AesSbox.scala 41:63]
  wire  _T_3480 = _T_3478 ^ _T_3476; // @[AesSbox.scala 40:63]
  wire  _T_3482 = _T_3398 & _T_3415; // @[AesSbox.scala 41:63]
  wire  _T_3484 = _T_3482 ^ _T_3476; // @[AesSbox.scala 40:63]
  wire  _T_3486 = _T_3460 ^ _T_3458; // @[AesSbox.scala 40:63]
  wire  _T_3488 = _T_3464 ^ _T_3403; // @[AesSbox.scala 40:63]
  wire  _T_3490 = _T_3470 ^ _T_3468; // @[AesSbox.scala 40:63]
  wire  _T_3492 = _T_3474 ^ _T_3484; // @[AesSbox.scala 40:63]
  wire  _T_3494 = _T_3486 ^ _T_3480; // @[AesSbox.scala 40:63]
  wire  _T_3496 = _T_3488 ^ _T_3484; // @[AesSbox.scala 40:63]
  wire  _T_3498 = _T_3490 ^ _T_3480; // @[AesSbox.scala 40:63]
  wire  _T_3500 = _T_3492 ^ _T_3422; // @[AesSbox.scala 40:63]
  wire  _T_3502 = _T_3498 ^ _T_3500; // @[AesSbox.scala 40:63]
  wire  _T_3504 = _T_3498 & _T_3494; // @[AesSbox.scala 41:63]
  wire  _T_3506 = _T_3496 ^ _T_3504; // @[AesSbox.scala 40:63]
  wire  _T_3508 = _T_3494 ^ _T_3496; // @[AesSbox.scala 40:63]
  wire  _T_3510 = _T_3500 ^ _T_3504; // @[AesSbox.scala 40:63]
  wire  _T_3512 = _T_3510 & _T_3508; // @[AesSbox.scala 41:63]
  wire  _T_3514 = _T_3506 & _T_3502; // @[AesSbox.scala 41:63]
  wire  _T_3516 = _T_3494 & _T_3500; // @[AesSbox.scala 41:63]
  wire  _T_3518 = _T_3508 & _T_3516; // @[AesSbox.scala 41:63]
  wire  _T_3520 = _T_3508 ^ _T_3504; // @[AesSbox.scala 40:63]
  wire  _T_3522 = _T_3496 & _T_3498; // @[AesSbox.scala 41:63]
  wire  _T_3524 = _T_3502 & _T_3522; // @[AesSbox.scala 41:63]
  wire  _T_3526 = _T_3502 ^ _T_3504; // @[AesSbox.scala 40:63]
  wire  _T_3528 = _T_3496 ^ _T_3512; // @[AesSbox.scala 40:63]
  wire  _T_3530 = _T_3518 ^ _T_3520; // @[AesSbox.scala 40:63]
  wire  _T_3532 = _T_3500 ^ _T_3514; // @[AesSbox.scala 40:63]
  wire  _T_3534 = _T_3524 ^ _T_3526; // @[AesSbox.scala 40:63]
  wire  _T_3536 = _T_3530 ^ _T_3534; // @[AesSbox.scala 40:63]
  wire  _T_3538 = _T_3528 ^ _T_3532; // @[AesSbox.scala 40:63]
  wire  _T_3540 = _T_3528 ^ _T_3530; // @[AesSbox.scala 40:63]
  wire  _T_3542 = _T_3532 ^ _T_3534; // @[AesSbox.scala 40:63]
  wire  _T_3544 = _T_3538 ^ _T_3536; // @[AesSbox.scala 40:63]
  wire  _T_3546 = _T_3542 & _T_3444; // @[AesSbox.scala 41:63]
  wire  _T_3548 = _T_3534 & _T_3408; // @[AesSbox.scala 41:63]
  wire  _T_3550 = _T_3532 & _T_3442; // @[AesSbox.scala 41:63]
  wire  _T_3552 = _T_3540 & _T_3446; // @[AesSbox.scala 41:63]
  wire  _T_3554 = _T_3530 & _T_3413; // @[AesSbox.scala 41:63]
  wire  _T_3556 = _T_3528 & _T_3427; // @[AesSbox.scala 41:63]
  wire  _T_3558 = _T_3538 & _T_3450; // @[AesSbox.scala 41:63]
  wire  _T_3560 = _T_3544 & _T_3448; // @[AesSbox.scala 41:63]
  wire  _T_3562 = _T_3536 & _T_3415; // @[AesSbox.scala 41:63]
  wire  _T_3564 = _T_3542 & _T_3417; // @[AesSbox.scala 41:63]
  wire  _T_3566 = _T_3534 & _T_3392; // @[AesSbox.scala 41:63]
  wire  _T_3568 = _T_3532 & _T_3410; // @[AesSbox.scala 41:63]
  wire  _T_3570 = _T_3540 & _T_3419; // @[AesSbox.scala 41:63]
  wire  _T_3572 = _T_3530 & _T_3395; // @[AesSbox.scala 41:63]
  wire  _T_3574 = _T_3528 & _T_3429; // @[AesSbox.scala 41:63]
  wire  _T_3576 = _T_3538 & _T_3400; // @[AesSbox.scala 41:63]
  wire  _T_3578 = _T_3544 & _T_3431; // @[AesSbox.scala 41:63]
  wire  _T_3580 = _T_3536 & _T_3398; // @[AesSbox.scala 41:63]
  wire  _T_3582 = _T_3558 ^ _T_3576; // @[AesSbox.scala 40:63]
  wire  _T_3584 = _T_3570 ^ _T_3572; // @[AesSbox.scala 40:63]
  wire  _T_3586 = _T_3562 ^ _T_3578; // @[AesSbox.scala 40:63]
  wire  _T_3588 = _T_3548 ^ _T_3554; // @[AesSbox.scala 40:63]
  wire  _T_3590 = _T_3550 ^ _T_3566; // @[AesSbox.scala 40:63]
  wire  _T_3592 = _T_3546 ^ _T_3556; // @[AesSbox.scala 40:63]
  wire  _T_3594 = _T_3552 ^ _T_3574; // @[AesSbox.scala 40:63]
  wire  _T_3596 = _T_3582 ^ _T_3584; // @[AesSbox.scala 40:63]
  wire  _T_3598 = _T_3554 ^ _T_3560; // @[AesSbox.scala 40:63]
  wire  _T_3600 = _T_3564 ^ _T_3580; // @[AesSbox.scala 40:63]
  wire  _T_3602 = _T_3568 ^ _T_3590; // @[AesSbox.scala 40:63]
  wire  _T_3604 = _T_3582 ^ _T_3588; // @[AesSbox.scala 40:63]
  wire  _T_3606 = _T_3546 ^ _T_3550; // @[AesSbox.scala 40:63]
  wire  _T_3608 = _T_3552 ^ _T_3556; // @[AesSbox.scala 40:63]
  wire  _T_3610 = _T_3552 ^ _T_3578; // @[AesSbox.scala 40:63]
  wire  _T_3612 = _T_3562 ^ _T_3572; // @[AesSbox.scala 40:63]
  wire  _T_3614 = _T_3568 ^ _T_3576; // @[AesSbox.scala 40:63]
  wire  _T_3616 = _T_3570 ^ _T_3586; // @[AesSbox.scala 40:63]
  wire  _T_3618 = _T_3580 ^ _T_3592; // @[AesSbox.scala 40:63]
  wire  _T_3620 = _T_3586 ^ _T_3588; // @[AesSbox.scala 40:63]
  wire  _T_3622 = _T_3590 ^ _T_3594; // @[AesSbox.scala 40:63]
  wire  _T_3624 = _T_3586 ^ _T_3596; // @[AesSbox.scala 40:63]
  wire  _T_3626 = _T_3596 ^ _T_3598; // @[AesSbox.scala 40:63]
  wire  _T_3628 = _T_3592 ^ _T_3596; // @[AesSbox.scala 40:63]
  wire  _T_3630 = _T_3594 ^ _T_3602; // @[AesSbox.scala 40:63]
  wire  _T_3632 = _T_3600 ^ _T_3604; // @[AesSbox.scala 40:63]
  wire  _T_3634 = _T_3602 ^ _T_3618; // @[AesSbox.scala 40:63]
  wire  _T_3636 = _T_3604 ^ _T_3630; // @[AesSbox.scala 40:63]
  wire  _T_3638 = _T_3612 ^ _T_3622; // @[AesSbox.scala 40:63]
  wire  _T_3639 = _T_3608 ^ _T_3624; // @[AesSbox.scala 40:63]
  wire  _T_3640 = _T_3632 ^ _T_3638; // @[AesSbox.scala 40:63]
  wire  _T_3641 = _T_3616 ^ _T_3636; // @[AesSbox.scala 40:63]
  wire  _T_3642 = _T_3606 ^ _T_3624; // @[AesSbox.scala 40:63]
  wire  _T_3643 = _T_3626 ^ _T_3634; // @[AesSbox.scala 40:63]
  wire  _T_3644 = _T_3620 ^ _T_3628; // @[AesSbox.scala 40:63]
  wire  _T_3645 = _T_3610 ^ _T_3626; // @[AesSbox.scala 40:63]
  wire  _T_3646 = _T_3600 ^ _T_3614; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_3_0 = {_T_3639,_T_3640,_T_3641,_T_3642,_T_3643,_T_3644,_T_3645,_T_3646}; // @[Cat.scala 29:58]
  wire  _T_3671 = matrix_2_1[7] ^ matrix_2_1[4]; // @[AesSbox.scala 40:63]
  wire  _T_3673 = matrix_2_1[6] ^ matrix_2_1[4]; // @[AesSbox.scala 42:65]
  wire  _T_3674 = ~_T_3673; // @[AesSbox.scala 42:51]
  wire  _T_3676 = matrix_2_1[7] ^ matrix_2_1[6]; // @[AesSbox.scala 42:65]
  wire  _T_3677 = ~_T_3676; // @[AesSbox.scala 42:51]
  wire  _T_3679 = matrix_2_1[4] ^ matrix_2_1[3]; // @[AesSbox.scala 40:63]
  wire  _T_3681 = matrix_2_1[3] ^ matrix_2_1[0]; // @[AesSbox.scala 42:65]
  wire  _T_3682 = ~_T_3681; // @[AesSbox.scala 42:51]
  wire  _T_3684 = matrix_2_1[1] ^ matrix_2_1[0]; // @[AesSbox.scala 40:63]
  wire  _T_3686 = matrix_2_1[6] ^ _T_3671; // @[AesSbox.scala 42:65]
  wire  _T_3687 = ~_T_3686; // @[AesSbox.scala 42:51]
  wire  _T_3689 = _T_3674 ^ _T_3684; // @[AesSbox.scala 40:63]
  wire  _T_3691 = matrix_2_1[0] ^ _T_3679; // @[AesSbox.scala 42:65]
  wire  _T_3692 = ~_T_3691; // @[AesSbox.scala 42:51]
  wire  _T_3694 = _T_3677 ^ _T_3682; // @[AesSbox.scala 40:63]
  wire  _T_3696 = _T_3677 ^ _T_3684; // @[AesSbox.scala 40:63]
  wire  _T_3698 = _T_3679 ^ _T_3684; // @[AesSbox.scala 40:63]
  wire  _T_3700 = matrix_2_1[5] ^ _T_3679; // @[AesSbox.scala 42:65]
  wire  _T_3701 = ~_T_3700; // @[AesSbox.scala 42:51]
  wire  _T_3703 = matrix_2_1[6] ^ matrix_2_1[1]; // @[AesSbox.scala 40:63]
  wire  _T_3705 = matrix_2_1[5] ^ _T_3689; // @[AesSbox.scala 42:65]
  wire  _T_3706 = ~_T_3705; // @[AesSbox.scala 42:51]
  wire  _T_3708 = _T_3682 ^ _T_3703; // @[AesSbox.scala 40:63]
  wire  _T_3710 = matrix_2_1[3] ^ _T_3687; // @[AesSbox.scala 40:63]
  wire  _T_3712 = matrix_2_1[5] ^ matrix_2_1[2]; // @[AesSbox.scala 42:65]
  wire  _T_3713 = ~_T_3712; // @[AesSbox.scala 42:51]
  wire  _T_3715 = matrix_2_1[2] ^ matrix_2_1[1]; // @[AesSbox.scala 42:65]
  wire  _T_3716 = ~_T_3715; // @[AesSbox.scala 42:51]
  wire  _T_3718 = matrix_2_1[5] ^ matrix_2_1[3]; // @[AesSbox.scala 42:65]
  wire  _T_3719 = ~_T_3718; // @[AesSbox.scala 42:51]
  wire  _T_3721 = matrix_2_1[7] ^ _T_3713; // @[AesSbox.scala 40:63]
  wire  _T_3723 = _T_3674 ^ _T_3713; // @[AesSbox.scala 40:63]
  wire  _T_3725 = _T_3703 ^ _T_3719; // @[AesSbox.scala 40:63]
  wire  _T_3727 = _T_3679 ^ _T_3716; // @[AesSbox.scala 40:63]
  wire  _T_3729 = _T_3694 ^ _T_3727; // @[AesSbox.scala 40:63]
  wire  _T_3731 = _T_3694 ^ _T_3716; // @[AesSbox.scala 40:63]
  wire  _T_3733 = _T_3698 ^ _T_3725; // @[AesSbox.scala 40:63]
  wire  _T_3735 = _T_3696 & _T_3723; // @[AesSbox.scala 41:63]
  wire  _T_3737 = _T_3671 & _T_3687; // @[AesSbox.scala 41:63]
  wire  _T_3739 = _T_3731 ^ _T_3735; // @[AesSbox.scala 40:63]
  wire  _T_3741 = _T_3689 & _T_3721; // @[AesSbox.scala 41:63]
  wire  _T_3743 = _T_3741 ^ _T_3735; // @[AesSbox.scala 40:63]
  wire  _T_3745 = _T_3698 & _T_3725; // @[AesSbox.scala 41:63]
  wire  _T_3747 = _T_3674 & _T_3692; // @[AesSbox.scala 41:63]
  wire  _T_3749 = _T_3733 ^ _T_3745; // @[AesSbox.scala 40:63]
  wire  _T_3751 = _T_3708 & _T_3706; // @[AesSbox.scala 41:63]
  wire  _T_3753 = _T_3751 ^ _T_3745; // @[AesSbox.scala 40:63]
  wire  _T_3755 = _T_3679 & _T_3729; // @[AesSbox.scala 41:63]
  wire  _T_3757 = _T_3710 & _T_3727; // @[AesSbox.scala 41:63]
  wire  _T_3759 = _T_3757 ^ _T_3755; // @[AesSbox.scala 40:63]
  wire  _T_3761 = _T_3677 & _T_3694; // @[AesSbox.scala 41:63]
  wire  _T_3763 = _T_3761 ^ _T_3755; // @[AesSbox.scala 40:63]
  wire  _T_3765 = _T_3739 ^ _T_3737; // @[AesSbox.scala 40:63]
  wire  _T_3767 = _T_3743 ^ _T_3682; // @[AesSbox.scala 40:63]
  wire  _T_3769 = _T_3749 ^ _T_3747; // @[AesSbox.scala 40:63]
  wire  _T_3771 = _T_3753 ^ _T_3763; // @[AesSbox.scala 40:63]
  wire  _T_3773 = _T_3765 ^ _T_3759; // @[AesSbox.scala 40:63]
  wire  _T_3775 = _T_3767 ^ _T_3763; // @[AesSbox.scala 40:63]
  wire  _T_3777 = _T_3769 ^ _T_3759; // @[AesSbox.scala 40:63]
  wire  _T_3779 = _T_3771 ^ _T_3701; // @[AesSbox.scala 40:63]
  wire  _T_3781 = _T_3777 ^ _T_3779; // @[AesSbox.scala 40:63]
  wire  _T_3783 = _T_3777 & _T_3773; // @[AesSbox.scala 41:63]
  wire  _T_3785 = _T_3775 ^ _T_3783; // @[AesSbox.scala 40:63]
  wire  _T_3787 = _T_3773 ^ _T_3775; // @[AesSbox.scala 40:63]
  wire  _T_3789 = _T_3779 ^ _T_3783; // @[AesSbox.scala 40:63]
  wire  _T_3791 = _T_3789 & _T_3787; // @[AesSbox.scala 41:63]
  wire  _T_3793 = _T_3785 & _T_3781; // @[AesSbox.scala 41:63]
  wire  _T_3795 = _T_3773 & _T_3779; // @[AesSbox.scala 41:63]
  wire  _T_3797 = _T_3787 & _T_3795; // @[AesSbox.scala 41:63]
  wire  _T_3799 = _T_3787 ^ _T_3783; // @[AesSbox.scala 40:63]
  wire  _T_3801 = _T_3775 & _T_3777; // @[AesSbox.scala 41:63]
  wire  _T_3803 = _T_3781 & _T_3801; // @[AesSbox.scala 41:63]
  wire  _T_3805 = _T_3781 ^ _T_3783; // @[AesSbox.scala 40:63]
  wire  _T_3807 = _T_3775 ^ _T_3791; // @[AesSbox.scala 40:63]
  wire  _T_3809 = _T_3797 ^ _T_3799; // @[AesSbox.scala 40:63]
  wire  _T_3811 = _T_3779 ^ _T_3793; // @[AesSbox.scala 40:63]
  wire  _T_3813 = _T_3803 ^ _T_3805; // @[AesSbox.scala 40:63]
  wire  _T_3815 = _T_3809 ^ _T_3813; // @[AesSbox.scala 40:63]
  wire  _T_3817 = _T_3807 ^ _T_3811; // @[AesSbox.scala 40:63]
  wire  _T_3819 = _T_3807 ^ _T_3809; // @[AesSbox.scala 40:63]
  wire  _T_3821 = _T_3811 ^ _T_3813; // @[AesSbox.scala 40:63]
  wire  _T_3823 = _T_3817 ^ _T_3815; // @[AesSbox.scala 40:63]
  wire  _T_3825 = _T_3821 & _T_3723; // @[AesSbox.scala 41:63]
  wire  _T_3827 = _T_3813 & _T_3687; // @[AesSbox.scala 41:63]
  wire  _T_3829 = _T_3811 & _T_3721; // @[AesSbox.scala 41:63]
  wire  _T_3831 = _T_3819 & _T_3725; // @[AesSbox.scala 41:63]
  wire  _T_3833 = _T_3809 & _T_3692; // @[AesSbox.scala 41:63]
  wire  _T_3835 = _T_3807 & _T_3706; // @[AesSbox.scala 41:63]
  wire  _T_3837 = _T_3817 & _T_3729; // @[AesSbox.scala 41:63]
  wire  _T_3839 = _T_3823 & _T_3727; // @[AesSbox.scala 41:63]
  wire  _T_3841 = _T_3815 & _T_3694; // @[AesSbox.scala 41:63]
  wire  _T_3843 = _T_3821 & _T_3696; // @[AesSbox.scala 41:63]
  wire  _T_3845 = _T_3813 & _T_3671; // @[AesSbox.scala 41:63]
  wire  _T_3847 = _T_3811 & _T_3689; // @[AesSbox.scala 41:63]
  wire  _T_3849 = _T_3819 & _T_3698; // @[AesSbox.scala 41:63]
  wire  _T_3851 = _T_3809 & _T_3674; // @[AesSbox.scala 41:63]
  wire  _T_3853 = _T_3807 & _T_3708; // @[AesSbox.scala 41:63]
  wire  _T_3855 = _T_3817 & _T_3679; // @[AesSbox.scala 41:63]
  wire  _T_3857 = _T_3823 & _T_3710; // @[AesSbox.scala 41:63]
  wire  _T_3859 = _T_3815 & _T_3677; // @[AesSbox.scala 41:63]
  wire  _T_3861 = _T_3837 ^ _T_3855; // @[AesSbox.scala 40:63]
  wire  _T_3863 = _T_3849 ^ _T_3851; // @[AesSbox.scala 40:63]
  wire  _T_3865 = _T_3841 ^ _T_3857; // @[AesSbox.scala 40:63]
  wire  _T_3867 = _T_3827 ^ _T_3833; // @[AesSbox.scala 40:63]
  wire  _T_3869 = _T_3829 ^ _T_3845; // @[AesSbox.scala 40:63]
  wire  _T_3871 = _T_3825 ^ _T_3835; // @[AesSbox.scala 40:63]
  wire  _T_3873 = _T_3831 ^ _T_3853; // @[AesSbox.scala 40:63]
  wire  _T_3875 = _T_3861 ^ _T_3863; // @[AesSbox.scala 40:63]
  wire  _T_3877 = _T_3833 ^ _T_3839; // @[AesSbox.scala 40:63]
  wire  _T_3879 = _T_3843 ^ _T_3859; // @[AesSbox.scala 40:63]
  wire  _T_3881 = _T_3847 ^ _T_3869; // @[AesSbox.scala 40:63]
  wire  _T_3883 = _T_3861 ^ _T_3867; // @[AesSbox.scala 40:63]
  wire  _T_3885 = _T_3825 ^ _T_3829; // @[AesSbox.scala 40:63]
  wire  _T_3887 = _T_3831 ^ _T_3835; // @[AesSbox.scala 40:63]
  wire  _T_3889 = _T_3831 ^ _T_3857; // @[AesSbox.scala 40:63]
  wire  _T_3891 = _T_3841 ^ _T_3851; // @[AesSbox.scala 40:63]
  wire  _T_3893 = _T_3847 ^ _T_3855; // @[AesSbox.scala 40:63]
  wire  _T_3895 = _T_3849 ^ _T_3865; // @[AesSbox.scala 40:63]
  wire  _T_3897 = _T_3859 ^ _T_3871; // @[AesSbox.scala 40:63]
  wire  _T_3899 = _T_3865 ^ _T_3867; // @[AesSbox.scala 40:63]
  wire  _T_3901 = _T_3869 ^ _T_3873; // @[AesSbox.scala 40:63]
  wire  _T_3903 = _T_3865 ^ _T_3875; // @[AesSbox.scala 40:63]
  wire  _T_3905 = _T_3875 ^ _T_3877; // @[AesSbox.scala 40:63]
  wire  _T_3907 = _T_3871 ^ _T_3875; // @[AesSbox.scala 40:63]
  wire  _T_3909 = _T_3873 ^ _T_3881; // @[AesSbox.scala 40:63]
  wire  _T_3911 = _T_3879 ^ _T_3883; // @[AesSbox.scala 40:63]
  wire  _T_3913 = _T_3881 ^ _T_3897; // @[AesSbox.scala 40:63]
  wire  _T_3915 = _T_3883 ^ _T_3909; // @[AesSbox.scala 40:63]
  wire  _T_3917 = _T_3891 ^ _T_3901; // @[AesSbox.scala 40:63]
  wire  _T_3918 = _T_3887 ^ _T_3903; // @[AesSbox.scala 40:63]
  wire  _T_3919 = _T_3911 ^ _T_3917; // @[AesSbox.scala 40:63]
  wire  _T_3920 = _T_3895 ^ _T_3915; // @[AesSbox.scala 40:63]
  wire  _T_3921 = _T_3885 ^ _T_3903; // @[AesSbox.scala 40:63]
  wire  _T_3922 = _T_3905 ^ _T_3913; // @[AesSbox.scala 40:63]
  wire  _T_3923 = _T_3899 ^ _T_3907; // @[AesSbox.scala 40:63]
  wire  _T_3924 = _T_3889 ^ _T_3905; // @[AesSbox.scala 40:63]
  wire  _T_3925 = _T_3879 ^ _T_3893; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_3_1 = {_T_3918,_T_3919,_T_3920,_T_3921,_T_3922,_T_3923,_T_3924,_T_3925}; // @[Cat.scala 29:58]
  wire  _T_3950 = matrix_1_2[7] ^ matrix_1_2[4]; // @[AesSbox.scala 40:63]
  wire  _T_3952 = matrix_1_2[6] ^ matrix_1_2[4]; // @[AesSbox.scala 42:65]
  wire  _T_3953 = ~_T_3952; // @[AesSbox.scala 42:51]
  wire  _T_3955 = matrix_1_2[7] ^ matrix_1_2[6]; // @[AesSbox.scala 42:65]
  wire  _T_3956 = ~_T_3955; // @[AesSbox.scala 42:51]
  wire  _T_3958 = matrix_1_2[4] ^ matrix_1_2[3]; // @[AesSbox.scala 40:63]
  wire  _T_3960 = matrix_1_2[3] ^ matrix_1_2[0]; // @[AesSbox.scala 42:65]
  wire  _T_3961 = ~_T_3960; // @[AesSbox.scala 42:51]
  wire  _T_3963 = matrix_1_2[1] ^ matrix_1_2[0]; // @[AesSbox.scala 40:63]
  wire  _T_3965 = matrix_1_2[6] ^ _T_3950; // @[AesSbox.scala 42:65]
  wire  _T_3966 = ~_T_3965; // @[AesSbox.scala 42:51]
  wire  _T_3968 = _T_3953 ^ _T_3963; // @[AesSbox.scala 40:63]
  wire  _T_3970 = matrix_1_2[0] ^ _T_3958; // @[AesSbox.scala 42:65]
  wire  _T_3971 = ~_T_3970; // @[AesSbox.scala 42:51]
  wire  _T_3973 = _T_3956 ^ _T_3961; // @[AesSbox.scala 40:63]
  wire  _T_3975 = _T_3956 ^ _T_3963; // @[AesSbox.scala 40:63]
  wire  _T_3977 = _T_3958 ^ _T_3963; // @[AesSbox.scala 40:63]
  wire  _T_3979 = matrix_1_2[5] ^ _T_3958; // @[AesSbox.scala 42:65]
  wire  _T_3980 = ~_T_3979; // @[AesSbox.scala 42:51]
  wire  _T_3982 = matrix_1_2[6] ^ matrix_1_2[1]; // @[AesSbox.scala 40:63]
  wire  _T_3984 = matrix_1_2[5] ^ _T_3968; // @[AesSbox.scala 42:65]
  wire  _T_3985 = ~_T_3984; // @[AesSbox.scala 42:51]
  wire  _T_3987 = _T_3961 ^ _T_3982; // @[AesSbox.scala 40:63]
  wire  _T_3989 = matrix_1_2[3] ^ _T_3966; // @[AesSbox.scala 40:63]
  wire  _T_3991 = matrix_1_2[5] ^ matrix_1_2[2]; // @[AesSbox.scala 42:65]
  wire  _T_3992 = ~_T_3991; // @[AesSbox.scala 42:51]
  wire  _T_3994 = matrix_1_2[2] ^ matrix_1_2[1]; // @[AesSbox.scala 42:65]
  wire  _T_3995 = ~_T_3994; // @[AesSbox.scala 42:51]
  wire  _T_3997 = matrix_1_2[5] ^ matrix_1_2[3]; // @[AesSbox.scala 42:65]
  wire  _T_3998 = ~_T_3997; // @[AesSbox.scala 42:51]
  wire  _T_4000 = matrix_1_2[7] ^ _T_3992; // @[AesSbox.scala 40:63]
  wire  _T_4002 = _T_3953 ^ _T_3992; // @[AesSbox.scala 40:63]
  wire  _T_4004 = _T_3982 ^ _T_3998; // @[AesSbox.scala 40:63]
  wire  _T_4006 = _T_3958 ^ _T_3995; // @[AesSbox.scala 40:63]
  wire  _T_4008 = _T_3973 ^ _T_4006; // @[AesSbox.scala 40:63]
  wire  _T_4010 = _T_3973 ^ _T_3995; // @[AesSbox.scala 40:63]
  wire  _T_4012 = _T_3977 ^ _T_4004; // @[AesSbox.scala 40:63]
  wire  _T_4014 = _T_3975 & _T_4002; // @[AesSbox.scala 41:63]
  wire  _T_4016 = _T_3950 & _T_3966; // @[AesSbox.scala 41:63]
  wire  _T_4018 = _T_4010 ^ _T_4014; // @[AesSbox.scala 40:63]
  wire  _T_4020 = _T_3968 & _T_4000; // @[AesSbox.scala 41:63]
  wire  _T_4022 = _T_4020 ^ _T_4014; // @[AesSbox.scala 40:63]
  wire  _T_4024 = _T_3977 & _T_4004; // @[AesSbox.scala 41:63]
  wire  _T_4026 = _T_3953 & _T_3971; // @[AesSbox.scala 41:63]
  wire  _T_4028 = _T_4012 ^ _T_4024; // @[AesSbox.scala 40:63]
  wire  _T_4030 = _T_3987 & _T_3985; // @[AesSbox.scala 41:63]
  wire  _T_4032 = _T_4030 ^ _T_4024; // @[AesSbox.scala 40:63]
  wire  _T_4034 = _T_3958 & _T_4008; // @[AesSbox.scala 41:63]
  wire  _T_4036 = _T_3989 & _T_4006; // @[AesSbox.scala 41:63]
  wire  _T_4038 = _T_4036 ^ _T_4034; // @[AesSbox.scala 40:63]
  wire  _T_4040 = _T_3956 & _T_3973; // @[AesSbox.scala 41:63]
  wire  _T_4042 = _T_4040 ^ _T_4034; // @[AesSbox.scala 40:63]
  wire  _T_4044 = _T_4018 ^ _T_4016; // @[AesSbox.scala 40:63]
  wire  _T_4046 = _T_4022 ^ _T_3961; // @[AesSbox.scala 40:63]
  wire  _T_4048 = _T_4028 ^ _T_4026; // @[AesSbox.scala 40:63]
  wire  _T_4050 = _T_4032 ^ _T_4042; // @[AesSbox.scala 40:63]
  wire  _T_4052 = _T_4044 ^ _T_4038; // @[AesSbox.scala 40:63]
  wire  _T_4054 = _T_4046 ^ _T_4042; // @[AesSbox.scala 40:63]
  wire  _T_4056 = _T_4048 ^ _T_4038; // @[AesSbox.scala 40:63]
  wire  _T_4058 = _T_4050 ^ _T_3980; // @[AesSbox.scala 40:63]
  wire  _T_4060 = _T_4056 ^ _T_4058; // @[AesSbox.scala 40:63]
  wire  _T_4062 = _T_4056 & _T_4052; // @[AesSbox.scala 41:63]
  wire  _T_4064 = _T_4054 ^ _T_4062; // @[AesSbox.scala 40:63]
  wire  _T_4066 = _T_4052 ^ _T_4054; // @[AesSbox.scala 40:63]
  wire  _T_4068 = _T_4058 ^ _T_4062; // @[AesSbox.scala 40:63]
  wire  _T_4070 = _T_4068 & _T_4066; // @[AesSbox.scala 41:63]
  wire  _T_4072 = _T_4064 & _T_4060; // @[AesSbox.scala 41:63]
  wire  _T_4074 = _T_4052 & _T_4058; // @[AesSbox.scala 41:63]
  wire  _T_4076 = _T_4066 & _T_4074; // @[AesSbox.scala 41:63]
  wire  _T_4078 = _T_4066 ^ _T_4062; // @[AesSbox.scala 40:63]
  wire  _T_4080 = _T_4054 & _T_4056; // @[AesSbox.scala 41:63]
  wire  _T_4082 = _T_4060 & _T_4080; // @[AesSbox.scala 41:63]
  wire  _T_4084 = _T_4060 ^ _T_4062; // @[AesSbox.scala 40:63]
  wire  _T_4086 = _T_4054 ^ _T_4070; // @[AesSbox.scala 40:63]
  wire  _T_4088 = _T_4076 ^ _T_4078; // @[AesSbox.scala 40:63]
  wire  _T_4090 = _T_4058 ^ _T_4072; // @[AesSbox.scala 40:63]
  wire  _T_4092 = _T_4082 ^ _T_4084; // @[AesSbox.scala 40:63]
  wire  _T_4094 = _T_4088 ^ _T_4092; // @[AesSbox.scala 40:63]
  wire  _T_4096 = _T_4086 ^ _T_4090; // @[AesSbox.scala 40:63]
  wire  _T_4098 = _T_4086 ^ _T_4088; // @[AesSbox.scala 40:63]
  wire  _T_4100 = _T_4090 ^ _T_4092; // @[AesSbox.scala 40:63]
  wire  _T_4102 = _T_4096 ^ _T_4094; // @[AesSbox.scala 40:63]
  wire  _T_4104 = _T_4100 & _T_4002; // @[AesSbox.scala 41:63]
  wire  _T_4106 = _T_4092 & _T_3966; // @[AesSbox.scala 41:63]
  wire  _T_4108 = _T_4090 & _T_4000; // @[AesSbox.scala 41:63]
  wire  _T_4110 = _T_4098 & _T_4004; // @[AesSbox.scala 41:63]
  wire  _T_4112 = _T_4088 & _T_3971; // @[AesSbox.scala 41:63]
  wire  _T_4114 = _T_4086 & _T_3985; // @[AesSbox.scala 41:63]
  wire  _T_4116 = _T_4096 & _T_4008; // @[AesSbox.scala 41:63]
  wire  _T_4118 = _T_4102 & _T_4006; // @[AesSbox.scala 41:63]
  wire  _T_4120 = _T_4094 & _T_3973; // @[AesSbox.scala 41:63]
  wire  _T_4122 = _T_4100 & _T_3975; // @[AesSbox.scala 41:63]
  wire  _T_4124 = _T_4092 & _T_3950; // @[AesSbox.scala 41:63]
  wire  _T_4126 = _T_4090 & _T_3968; // @[AesSbox.scala 41:63]
  wire  _T_4128 = _T_4098 & _T_3977; // @[AesSbox.scala 41:63]
  wire  _T_4130 = _T_4088 & _T_3953; // @[AesSbox.scala 41:63]
  wire  _T_4132 = _T_4086 & _T_3987; // @[AesSbox.scala 41:63]
  wire  _T_4134 = _T_4096 & _T_3958; // @[AesSbox.scala 41:63]
  wire  _T_4136 = _T_4102 & _T_3989; // @[AesSbox.scala 41:63]
  wire  _T_4138 = _T_4094 & _T_3956; // @[AesSbox.scala 41:63]
  wire  _T_4140 = _T_4116 ^ _T_4134; // @[AesSbox.scala 40:63]
  wire  _T_4142 = _T_4128 ^ _T_4130; // @[AesSbox.scala 40:63]
  wire  _T_4144 = _T_4120 ^ _T_4136; // @[AesSbox.scala 40:63]
  wire  _T_4146 = _T_4106 ^ _T_4112; // @[AesSbox.scala 40:63]
  wire  _T_4148 = _T_4108 ^ _T_4124; // @[AesSbox.scala 40:63]
  wire  _T_4150 = _T_4104 ^ _T_4114; // @[AesSbox.scala 40:63]
  wire  _T_4152 = _T_4110 ^ _T_4132; // @[AesSbox.scala 40:63]
  wire  _T_4154 = _T_4140 ^ _T_4142; // @[AesSbox.scala 40:63]
  wire  _T_4156 = _T_4112 ^ _T_4118; // @[AesSbox.scala 40:63]
  wire  _T_4158 = _T_4122 ^ _T_4138; // @[AesSbox.scala 40:63]
  wire  _T_4160 = _T_4126 ^ _T_4148; // @[AesSbox.scala 40:63]
  wire  _T_4162 = _T_4140 ^ _T_4146; // @[AesSbox.scala 40:63]
  wire  _T_4164 = _T_4104 ^ _T_4108; // @[AesSbox.scala 40:63]
  wire  _T_4166 = _T_4110 ^ _T_4114; // @[AesSbox.scala 40:63]
  wire  _T_4168 = _T_4110 ^ _T_4136; // @[AesSbox.scala 40:63]
  wire  _T_4170 = _T_4120 ^ _T_4130; // @[AesSbox.scala 40:63]
  wire  _T_4172 = _T_4126 ^ _T_4134; // @[AesSbox.scala 40:63]
  wire  _T_4174 = _T_4128 ^ _T_4144; // @[AesSbox.scala 40:63]
  wire  _T_4176 = _T_4138 ^ _T_4150; // @[AesSbox.scala 40:63]
  wire  _T_4178 = _T_4144 ^ _T_4146; // @[AesSbox.scala 40:63]
  wire  _T_4180 = _T_4148 ^ _T_4152; // @[AesSbox.scala 40:63]
  wire  _T_4182 = _T_4144 ^ _T_4154; // @[AesSbox.scala 40:63]
  wire  _T_4184 = _T_4154 ^ _T_4156; // @[AesSbox.scala 40:63]
  wire  _T_4186 = _T_4150 ^ _T_4154; // @[AesSbox.scala 40:63]
  wire  _T_4188 = _T_4152 ^ _T_4160; // @[AesSbox.scala 40:63]
  wire  _T_4190 = _T_4158 ^ _T_4162; // @[AesSbox.scala 40:63]
  wire  _T_4192 = _T_4160 ^ _T_4176; // @[AesSbox.scala 40:63]
  wire  _T_4194 = _T_4162 ^ _T_4188; // @[AesSbox.scala 40:63]
  wire  _T_4196 = _T_4170 ^ _T_4180; // @[AesSbox.scala 40:63]
  wire  _T_4197 = _T_4166 ^ _T_4182; // @[AesSbox.scala 40:63]
  wire  _T_4198 = _T_4190 ^ _T_4196; // @[AesSbox.scala 40:63]
  wire  _T_4199 = _T_4174 ^ _T_4194; // @[AesSbox.scala 40:63]
  wire  _T_4200 = _T_4164 ^ _T_4182; // @[AesSbox.scala 40:63]
  wire  _T_4201 = _T_4184 ^ _T_4192; // @[AesSbox.scala 40:63]
  wire  _T_4202 = _T_4178 ^ _T_4186; // @[AesSbox.scala 40:63]
  wire  _T_4203 = _T_4168 ^ _T_4184; // @[AesSbox.scala 40:63]
  wire  _T_4204 = _T_4158 ^ _T_4172; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_3_2 = {_T_4197,_T_4198,_T_4199,_T_4200,_T_4201,_T_4202,_T_4203,_T_4204}; // @[Cat.scala 29:58]
  wire  _T_4229 = matrix_0_3[7] ^ matrix_0_3[4]; // @[AesSbox.scala 40:63]
  wire  _T_4231 = matrix_0_3[6] ^ matrix_0_3[4]; // @[AesSbox.scala 42:65]
  wire  _T_4232 = ~_T_4231; // @[AesSbox.scala 42:51]
  wire  _T_4234 = matrix_0_3[7] ^ matrix_0_3[6]; // @[AesSbox.scala 42:65]
  wire  _T_4235 = ~_T_4234; // @[AesSbox.scala 42:51]
  wire  _T_4237 = matrix_0_3[4] ^ matrix_0_3[3]; // @[AesSbox.scala 40:63]
  wire  _T_4239 = matrix_0_3[3] ^ matrix_0_3[0]; // @[AesSbox.scala 42:65]
  wire  _T_4240 = ~_T_4239; // @[AesSbox.scala 42:51]
  wire  _T_4242 = matrix_0_3[1] ^ matrix_0_3[0]; // @[AesSbox.scala 40:63]
  wire  _T_4244 = matrix_0_3[6] ^ _T_4229; // @[AesSbox.scala 42:65]
  wire  _T_4245 = ~_T_4244; // @[AesSbox.scala 42:51]
  wire  _T_4247 = _T_4232 ^ _T_4242; // @[AesSbox.scala 40:63]
  wire  _T_4249 = matrix_0_3[0] ^ _T_4237; // @[AesSbox.scala 42:65]
  wire  _T_4250 = ~_T_4249; // @[AesSbox.scala 42:51]
  wire  _T_4252 = _T_4235 ^ _T_4240; // @[AesSbox.scala 40:63]
  wire  _T_4254 = _T_4235 ^ _T_4242; // @[AesSbox.scala 40:63]
  wire  _T_4256 = _T_4237 ^ _T_4242; // @[AesSbox.scala 40:63]
  wire  _T_4258 = matrix_0_3[5] ^ _T_4237; // @[AesSbox.scala 42:65]
  wire  _T_4259 = ~_T_4258; // @[AesSbox.scala 42:51]
  wire  _T_4261 = matrix_0_3[6] ^ matrix_0_3[1]; // @[AesSbox.scala 40:63]
  wire  _T_4263 = matrix_0_3[5] ^ _T_4247; // @[AesSbox.scala 42:65]
  wire  _T_4264 = ~_T_4263; // @[AesSbox.scala 42:51]
  wire  _T_4266 = _T_4240 ^ _T_4261; // @[AesSbox.scala 40:63]
  wire  _T_4268 = matrix_0_3[3] ^ _T_4245; // @[AesSbox.scala 40:63]
  wire  _T_4270 = matrix_0_3[5] ^ matrix_0_3[2]; // @[AesSbox.scala 42:65]
  wire  _T_4271 = ~_T_4270; // @[AesSbox.scala 42:51]
  wire  _T_4273 = matrix_0_3[2] ^ matrix_0_3[1]; // @[AesSbox.scala 42:65]
  wire  _T_4274 = ~_T_4273; // @[AesSbox.scala 42:51]
  wire  _T_4276 = matrix_0_3[5] ^ matrix_0_3[3]; // @[AesSbox.scala 42:65]
  wire  _T_4277 = ~_T_4276; // @[AesSbox.scala 42:51]
  wire  _T_4279 = matrix_0_3[7] ^ _T_4271; // @[AesSbox.scala 40:63]
  wire  _T_4281 = _T_4232 ^ _T_4271; // @[AesSbox.scala 40:63]
  wire  _T_4283 = _T_4261 ^ _T_4277; // @[AesSbox.scala 40:63]
  wire  _T_4285 = _T_4237 ^ _T_4274; // @[AesSbox.scala 40:63]
  wire  _T_4287 = _T_4252 ^ _T_4285; // @[AesSbox.scala 40:63]
  wire  _T_4289 = _T_4252 ^ _T_4274; // @[AesSbox.scala 40:63]
  wire  _T_4291 = _T_4256 ^ _T_4283; // @[AesSbox.scala 40:63]
  wire  _T_4293 = _T_4254 & _T_4281; // @[AesSbox.scala 41:63]
  wire  _T_4295 = _T_4229 & _T_4245; // @[AesSbox.scala 41:63]
  wire  _T_4297 = _T_4289 ^ _T_4293; // @[AesSbox.scala 40:63]
  wire  _T_4299 = _T_4247 & _T_4279; // @[AesSbox.scala 41:63]
  wire  _T_4301 = _T_4299 ^ _T_4293; // @[AesSbox.scala 40:63]
  wire  _T_4303 = _T_4256 & _T_4283; // @[AesSbox.scala 41:63]
  wire  _T_4305 = _T_4232 & _T_4250; // @[AesSbox.scala 41:63]
  wire  _T_4307 = _T_4291 ^ _T_4303; // @[AesSbox.scala 40:63]
  wire  _T_4309 = _T_4266 & _T_4264; // @[AesSbox.scala 41:63]
  wire  _T_4311 = _T_4309 ^ _T_4303; // @[AesSbox.scala 40:63]
  wire  _T_4313 = _T_4237 & _T_4287; // @[AesSbox.scala 41:63]
  wire  _T_4315 = _T_4268 & _T_4285; // @[AesSbox.scala 41:63]
  wire  _T_4317 = _T_4315 ^ _T_4313; // @[AesSbox.scala 40:63]
  wire  _T_4319 = _T_4235 & _T_4252; // @[AesSbox.scala 41:63]
  wire  _T_4321 = _T_4319 ^ _T_4313; // @[AesSbox.scala 40:63]
  wire  _T_4323 = _T_4297 ^ _T_4295; // @[AesSbox.scala 40:63]
  wire  _T_4325 = _T_4301 ^ _T_4240; // @[AesSbox.scala 40:63]
  wire  _T_4327 = _T_4307 ^ _T_4305; // @[AesSbox.scala 40:63]
  wire  _T_4329 = _T_4311 ^ _T_4321; // @[AesSbox.scala 40:63]
  wire  _T_4331 = _T_4323 ^ _T_4317; // @[AesSbox.scala 40:63]
  wire  _T_4333 = _T_4325 ^ _T_4321; // @[AesSbox.scala 40:63]
  wire  _T_4335 = _T_4327 ^ _T_4317; // @[AesSbox.scala 40:63]
  wire  _T_4337 = _T_4329 ^ _T_4259; // @[AesSbox.scala 40:63]
  wire  _T_4339 = _T_4335 ^ _T_4337; // @[AesSbox.scala 40:63]
  wire  _T_4341 = _T_4335 & _T_4331; // @[AesSbox.scala 41:63]
  wire  _T_4343 = _T_4333 ^ _T_4341; // @[AesSbox.scala 40:63]
  wire  _T_4345 = _T_4331 ^ _T_4333; // @[AesSbox.scala 40:63]
  wire  _T_4347 = _T_4337 ^ _T_4341; // @[AesSbox.scala 40:63]
  wire  _T_4349 = _T_4347 & _T_4345; // @[AesSbox.scala 41:63]
  wire  _T_4351 = _T_4343 & _T_4339; // @[AesSbox.scala 41:63]
  wire  _T_4353 = _T_4331 & _T_4337; // @[AesSbox.scala 41:63]
  wire  _T_4355 = _T_4345 & _T_4353; // @[AesSbox.scala 41:63]
  wire  _T_4357 = _T_4345 ^ _T_4341; // @[AesSbox.scala 40:63]
  wire  _T_4359 = _T_4333 & _T_4335; // @[AesSbox.scala 41:63]
  wire  _T_4361 = _T_4339 & _T_4359; // @[AesSbox.scala 41:63]
  wire  _T_4363 = _T_4339 ^ _T_4341; // @[AesSbox.scala 40:63]
  wire  _T_4365 = _T_4333 ^ _T_4349; // @[AesSbox.scala 40:63]
  wire  _T_4367 = _T_4355 ^ _T_4357; // @[AesSbox.scala 40:63]
  wire  _T_4369 = _T_4337 ^ _T_4351; // @[AesSbox.scala 40:63]
  wire  _T_4371 = _T_4361 ^ _T_4363; // @[AesSbox.scala 40:63]
  wire  _T_4373 = _T_4367 ^ _T_4371; // @[AesSbox.scala 40:63]
  wire  _T_4375 = _T_4365 ^ _T_4369; // @[AesSbox.scala 40:63]
  wire  _T_4377 = _T_4365 ^ _T_4367; // @[AesSbox.scala 40:63]
  wire  _T_4379 = _T_4369 ^ _T_4371; // @[AesSbox.scala 40:63]
  wire  _T_4381 = _T_4375 ^ _T_4373; // @[AesSbox.scala 40:63]
  wire  _T_4383 = _T_4379 & _T_4281; // @[AesSbox.scala 41:63]
  wire  _T_4385 = _T_4371 & _T_4245; // @[AesSbox.scala 41:63]
  wire  _T_4387 = _T_4369 & _T_4279; // @[AesSbox.scala 41:63]
  wire  _T_4389 = _T_4377 & _T_4283; // @[AesSbox.scala 41:63]
  wire  _T_4391 = _T_4367 & _T_4250; // @[AesSbox.scala 41:63]
  wire  _T_4393 = _T_4365 & _T_4264; // @[AesSbox.scala 41:63]
  wire  _T_4395 = _T_4375 & _T_4287; // @[AesSbox.scala 41:63]
  wire  _T_4397 = _T_4381 & _T_4285; // @[AesSbox.scala 41:63]
  wire  _T_4399 = _T_4373 & _T_4252; // @[AesSbox.scala 41:63]
  wire  _T_4401 = _T_4379 & _T_4254; // @[AesSbox.scala 41:63]
  wire  _T_4403 = _T_4371 & _T_4229; // @[AesSbox.scala 41:63]
  wire  _T_4405 = _T_4369 & _T_4247; // @[AesSbox.scala 41:63]
  wire  _T_4407 = _T_4377 & _T_4256; // @[AesSbox.scala 41:63]
  wire  _T_4409 = _T_4367 & _T_4232; // @[AesSbox.scala 41:63]
  wire  _T_4411 = _T_4365 & _T_4266; // @[AesSbox.scala 41:63]
  wire  _T_4413 = _T_4375 & _T_4237; // @[AesSbox.scala 41:63]
  wire  _T_4415 = _T_4381 & _T_4268; // @[AesSbox.scala 41:63]
  wire  _T_4417 = _T_4373 & _T_4235; // @[AesSbox.scala 41:63]
  wire  _T_4419 = _T_4395 ^ _T_4413; // @[AesSbox.scala 40:63]
  wire  _T_4421 = _T_4407 ^ _T_4409; // @[AesSbox.scala 40:63]
  wire  _T_4423 = _T_4399 ^ _T_4415; // @[AesSbox.scala 40:63]
  wire  _T_4425 = _T_4385 ^ _T_4391; // @[AesSbox.scala 40:63]
  wire  _T_4427 = _T_4387 ^ _T_4403; // @[AesSbox.scala 40:63]
  wire  _T_4429 = _T_4383 ^ _T_4393; // @[AesSbox.scala 40:63]
  wire  _T_4431 = _T_4389 ^ _T_4411; // @[AesSbox.scala 40:63]
  wire  _T_4433 = _T_4419 ^ _T_4421; // @[AesSbox.scala 40:63]
  wire  _T_4435 = _T_4391 ^ _T_4397; // @[AesSbox.scala 40:63]
  wire  _T_4437 = _T_4401 ^ _T_4417; // @[AesSbox.scala 40:63]
  wire  _T_4439 = _T_4405 ^ _T_4427; // @[AesSbox.scala 40:63]
  wire  _T_4441 = _T_4419 ^ _T_4425; // @[AesSbox.scala 40:63]
  wire  _T_4443 = _T_4383 ^ _T_4387; // @[AesSbox.scala 40:63]
  wire  _T_4445 = _T_4389 ^ _T_4393; // @[AesSbox.scala 40:63]
  wire  _T_4447 = _T_4389 ^ _T_4415; // @[AesSbox.scala 40:63]
  wire  _T_4449 = _T_4399 ^ _T_4409; // @[AesSbox.scala 40:63]
  wire  _T_4451 = _T_4405 ^ _T_4413; // @[AesSbox.scala 40:63]
  wire  _T_4453 = _T_4407 ^ _T_4423; // @[AesSbox.scala 40:63]
  wire  _T_4455 = _T_4417 ^ _T_4429; // @[AesSbox.scala 40:63]
  wire  _T_4457 = _T_4423 ^ _T_4425; // @[AesSbox.scala 40:63]
  wire  _T_4459 = _T_4427 ^ _T_4431; // @[AesSbox.scala 40:63]
  wire  _T_4461 = _T_4423 ^ _T_4433; // @[AesSbox.scala 40:63]
  wire  _T_4463 = _T_4433 ^ _T_4435; // @[AesSbox.scala 40:63]
  wire  _T_4465 = _T_4429 ^ _T_4433; // @[AesSbox.scala 40:63]
  wire  _T_4467 = _T_4431 ^ _T_4439; // @[AesSbox.scala 40:63]
  wire  _T_4469 = _T_4437 ^ _T_4441; // @[AesSbox.scala 40:63]
  wire  _T_4471 = _T_4439 ^ _T_4455; // @[AesSbox.scala 40:63]
  wire  _T_4473 = _T_4441 ^ _T_4467; // @[AesSbox.scala 40:63]
  wire  _T_4475 = _T_4449 ^ _T_4459; // @[AesSbox.scala 40:63]
  wire  _T_4476 = _T_4445 ^ _T_4461; // @[AesSbox.scala 40:63]
  wire  _T_4477 = _T_4469 ^ _T_4475; // @[AesSbox.scala 40:63]
  wire  _T_4478 = _T_4453 ^ _T_4473; // @[AesSbox.scala 40:63]
  wire  _T_4479 = _T_4443 ^ _T_4461; // @[AesSbox.scala 40:63]
  wire  _T_4480 = _T_4463 ^ _T_4471; // @[AesSbox.scala 40:63]
  wire  _T_4481 = _T_4457 ^ _T_4465; // @[AesSbox.scala 40:63]
  wire  _T_4482 = _T_4447 ^ _T_4463; // @[AesSbox.scala 40:63]
  wire  _T_4483 = _T_4437 ^ _T_4451; // @[AesSbox.scala 40:63]
  wire [7:0] roundPart1_3_3 = {_T_4476,_T_4477,_T_4478,_T_4479,_T_4480,_T_4481,_T_4482,_T_4483}; // @[Cat.scala 29:58]
  wire [3:0] keyEndAddr = io_aes256 ? 4'he : 4'ha; // @[AesDecrypt.scala 73:25]
  wire [7:0] _GEN_16 = 4'h1 == keyEndAddr ? io_keys_1_0_0 : io_keys_0_0_0; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_17 = 4'h1 == keyEndAddr ? io_keys_1_0_1 : io_keys_0_0_1; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_18 = 4'h1 == keyEndAddr ? io_keys_1_0_2 : io_keys_0_0_2; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_19 = 4'h1 == keyEndAddr ? io_keys_1_0_3 : io_keys_0_0_3; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_20 = 4'h1 == keyEndAddr ? io_keys_1_1_0 : io_keys_0_1_0; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_21 = 4'h1 == keyEndAddr ? io_keys_1_1_1 : io_keys_0_1_1; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_22 = 4'h1 == keyEndAddr ? io_keys_1_1_2 : io_keys_0_1_2; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_23 = 4'h1 == keyEndAddr ? io_keys_1_1_3 : io_keys_0_1_3; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_24 = 4'h1 == keyEndAddr ? io_keys_1_2_0 : io_keys_0_2_0; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_25 = 4'h1 == keyEndAddr ? io_keys_1_2_1 : io_keys_0_2_1; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_26 = 4'h1 == keyEndAddr ? io_keys_1_2_2 : io_keys_0_2_2; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_27 = 4'h1 == keyEndAddr ? io_keys_1_2_3 : io_keys_0_2_3; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_28 = 4'h1 == keyEndAddr ? io_keys_1_3_0 : io_keys_0_3_0; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_29 = 4'h1 == keyEndAddr ? io_keys_1_3_1 : io_keys_0_3_1; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_30 = 4'h1 == keyEndAddr ? io_keys_1_3_2 : io_keys_0_3_2; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_31 = 4'h1 == keyEndAddr ? io_keys_1_3_3 : io_keys_0_3_3; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_32 = 4'h2 == keyEndAddr ? io_keys_2_0_0 : _GEN_16; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_33 = 4'h2 == keyEndAddr ? io_keys_2_0_1 : _GEN_17; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_34 = 4'h2 == keyEndAddr ? io_keys_2_0_2 : _GEN_18; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_35 = 4'h2 == keyEndAddr ? io_keys_2_0_3 : _GEN_19; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_36 = 4'h2 == keyEndAddr ? io_keys_2_1_0 : _GEN_20; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_37 = 4'h2 == keyEndAddr ? io_keys_2_1_1 : _GEN_21; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_38 = 4'h2 == keyEndAddr ? io_keys_2_1_2 : _GEN_22; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_39 = 4'h2 == keyEndAddr ? io_keys_2_1_3 : _GEN_23; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_40 = 4'h2 == keyEndAddr ? io_keys_2_2_0 : _GEN_24; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_41 = 4'h2 == keyEndAddr ? io_keys_2_2_1 : _GEN_25; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_42 = 4'h2 == keyEndAddr ? io_keys_2_2_2 : _GEN_26; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_43 = 4'h2 == keyEndAddr ? io_keys_2_2_3 : _GEN_27; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_44 = 4'h2 == keyEndAddr ? io_keys_2_3_0 : _GEN_28; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_45 = 4'h2 == keyEndAddr ? io_keys_2_3_1 : _GEN_29; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_46 = 4'h2 == keyEndAddr ? io_keys_2_3_2 : _GEN_30; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_47 = 4'h2 == keyEndAddr ? io_keys_2_3_3 : _GEN_31; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_48 = 4'h3 == keyEndAddr ? io_keys_3_0_0 : _GEN_32; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_49 = 4'h3 == keyEndAddr ? io_keys_3_0_1 : _GEN_33; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_50 = 4'h3 == keyEndAddr ? io_keys_3_0_2 : _GEN_34; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_51 = 4'h3 == keyEndAddr ? io_keys_3_0_3 : _GEN_35; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_52 = 4'h3 == keyEndAddr ? io_keys_3_1_0 : _GEN_36; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_53 = 4'h3 == keyEndAddr ? io_keys_3_1_1 : _GEN_37; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_54 = 4'h3 == keyEndAddr ? io_keys_3_1_2 : _GEN_38; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_55 = 4'h3 == keyEndAddr ? io_keys_3_1_3 : _GEN_39; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_56 = 4'h3 == keyEndAddr ? io_keys_3_2_0 : _GEN_40; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_57 = 4'h3 == keyEndAddr ? io_keys_3_2_1 : _GEN_41; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_58 = 4'h3 == keyEndAddr ? io_keys_3_2_2 : _GEN_42; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_59 = 4'h3 == keyEndAddr ? io_keys_3_2_3 : _GEN_43; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_60 = 4'h3 == keyEndAddr ? io_keys_3_3_0 : _GEN_44; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_61 = 4'h3 == keyEndAddr ? io_keys_3_3_1 : _GEN_45; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_62 = 4'h3 == keyEndAddr ? io_keys_3_3_2 : _GEN_46; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_63 = 4'h3 == keyEndAddr ? io_keys_3_3_3 : _GEN_47; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_64 = 4'h4 == keyEndAddr ? io_keys_4_0_0 : _GEN_48; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_65 = 4'h4 == keyEndAddr ? io_keys_4_0_1 : _GEN_49; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_66 = 4'h4 == keyEndAddr ? io_keys_4_0_2 : _GEN_50; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_67 = 4'h4 == keyEndAddr ? io_keys_4_0_3 : _GEN_51; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_68 = 4'h4 == keyEndAddr ? io_keys_4_1_0 : _GEN_52; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_69 = 4'h4 == keyEndAddr ? io_keys_4_1_1 : _GEN_53; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_70 = 4'h4 == keyEndAddr ? io_keys_4_1_2 : _GEN_54; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_71 = 4'h4 == keyEndAddr ? io_keys_4_1_3 : _GEN_55; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_72 = 4'h4 == keyEndAddr ? io_keys_4_2_0 : _GEN_56; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_73 = 4'h4 == keyEndAddr ? io_keys_4_2_1 : _GEN_57; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_74 = 4'h4 == keyEndAddr ? io_keys_4_2_2 : _GEN_58; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_75 = 4'h4 == keyEndAddr ? io_keys_4_2_3 : _GEN_59; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_76 = 4'h4 == keyEndAddr ? io_keys_4_3_0 : _GEN_60; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_77 = 4'h4 == keyEndAddr ? io_keys_4_3_1 : _GEN_61; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_78 = 4'h4 == keyEndAddr ? io_keys_4_3_2 : _GEN_62; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_79 = 4'h4 == keyEndAddr ? io_keys_4_3_3 : _GEN_63; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_80 = 4'h5 == keyEndAddr ? io_keys_5_0_0 : _GEN_64; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_81 = 4'h5 == keyEndAddr ? io_keys_5_0_1 : _GEN_65; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_82 = 4'h5 == keyEndAddr ? io_keys_5_0_2 : _GEN_66; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_83 = 4'h5 == keyEndAddr ? io_keys_5_0_3 : _GEN_67; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_84 = 4'h5 == keyEndAddr ? io_keys_5_1_0 : _GEN_68; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_85 = 4'h5 == keyEndAddr ? io_keys_5_1_1 : _GEN_69; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_86 = 4'h5 == keyEndAddr ? io_keys_5_1_2 : _GEN_70; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_87 = 4'h5 == keyEndAddr ? io_keys_5_1_3 : _GEN_71; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_88 = 4'h5 == keyEndAddr ? io_keys_5_2_0 : _GEN_72; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_89 = 4'h5 == keyEndAddr ? io_keys_5_2_1 : _GEN_73; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_90 = 4'h5 == keyEndAddr ? io_keys_5_2_2 : _GEN_74; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_91 = 4'h5 == keyEndAddr ? io_keys_5_2_3 : _GEN_75; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_92 = 4'h5 == keyEndAddr ? io_keys_5_3_0 : _GEN_76; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_93 = 4'h5 == keyEndAddr ? io_keys_5_3_1 : _GEN_77; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_94 = 4'h5 == keyEndAddr ? io_keys_5_3_2 : _GEN_78; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_95 = 4'h5 == keyEndAddr ? io_keys_5_3_3 : _GEN_79; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_96 = 4'h6 == keyEndAddr ? io_keys_6_0_0 : _GEN_80; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_97 = 4'h6 == keyEndAddr ? io_keys_6_0_1 : _GEN_81; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_98 = 4'h6 == keyEndAddr ? io_keys_6_0_2 : _GEN_82; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_99 = 4'h6 == keyEndAddr ? io_keys_6_0_3 : _GEN_83; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_100 = 4'h6 == keyEndAddr ? io_keys_6_1_0 : _GEN_84; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_101 = 4'h6 == keyEndAddr ? io_keys_6_1_1 : _GEN_85; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_102 = 4'h6 == keyEndAddr ? io_keys_6_1_2 : _GEN_86; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_103 = 4'h6 == keyEndAddr ? io_keys_6_1_3 : _GEN_87; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_104 = 4'h6 == keyEndAddr ? io_keys_6_2_0 : _GEN_88; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_105 = 4'h6 == keyEndAddr ? io_keys_6_2_1 : _GEN_89; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_106 = 4'h6 == keyEndAddr ? io_keys_6_2_2 : _GEN_90; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_107 = 4'h6 == keyEndAddr ? io_keys_6_2_3 : _GEN_91; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_108 = 4'h6 == keyEndAddr ? io_keys_6_3_0 : _GEN_92; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_109 = 4'h6 == keyEndAddr ? io_keys_6_3_1 : _GEN_93; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_110 = 4'h6 == keyEndAddr ? io_keys_6_3_2 : _GEN_94; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_111 = 4'h6 == keyEndAddr ? io_keys_6_3_3 : _GEN_95; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_112 = 4'h7 == keyEndAddr ? io_keys_7_0_0 : _GEN_96; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_113 = 4'h7 == keyEndAddr ? io_keys_7_0_1 : _GEN_97; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_114 = 4'h7 == keyEndAddr ? io_keys_7_0_2 : _GEN_98; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_115 = 4'h7 == keyEndAddr ? io_keys_7_0_3 : _GEN_99; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_116 = 4'h7 == keyEndAddr ? io_keys_7_1_0 : _GEN_100; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_117 = 4'h7 == keyEndAddr ? io_keys_7_1_1 : _GEN_101; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_118 = 4'h7 == keyEndAddr ? io_keys_7_1_2 : _GEN_102; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_119 = 4'h7 == keyEndAddr ? io_keys_7_1_3 : _GEN_103; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_120 = 4'h7 == keyEndAddr ? io_keys_7_2_0 : _GEN_104; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_121 = 4'h7 == keyEndAddr ? io_keys_7_2_1 : _GEN_105; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_122 = 4'h7 == keyEndAddr ? io_keys_7_2_2 : _GEN_106; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_123 = 4'h7 == keyEndAddr ? io_keys_7_2_3 : _GEN_107; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_124 = 4'h7 == keyEndAddr ? io_keys_7_3_0 : _GEN_108; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_125 = 4'h7 == keyEndAddr ? io_keys_7_3_1 : _GEN_109; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_126 = 4'h7 == keyEndAddr ? io_keys_7_3_2 : _GEN_110; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_127 = 4'h7 == keyEndAddr ? io_keys_7_3_3 : _GEN_111; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_128 = 4'h8 == keyEndAddr ? io_keys_8_0_0 : _GEN_112; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_129 = 4'h8 == keyEndAddr ? io_keys_8_0_1 : _GEN_113; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_130 = 4'h8 == keyEndAddr ? io_keys_8_0_2 : _GEN_114; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_131 = 4'h8 == keyEndAddr ? io_keys_8_0_3 : _GEN_115; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_132 = 4'h8 == keyEndAddr ? io_keys_8_1_0 : _GEN_116; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_133 = 4'h8 == keyEndAddr ? io_keys_8_1_1 : _GEN_117; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_134 = 4'h8 == keyEndAddr ? io_keys_8_1_2 : _GEN_118; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_135 = 4'h8 == keyEndAddr ? io_keys_8_1_3 : _GEN_119; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_136 = 4'h8 == keyEndAddr ? io_keys_8_2_0 : _GEN_120; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_137 = 4'h8 == keyEndAddr ? io_keys_8_2_1 : _GEN_121; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_138 = 4'h8 == keyEndAddr ? io_keys_8_2_2 : _GEN_122; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_139 = 4'h8 == keyEndAddr ? io_keys_8_2_3 : _GEN_123; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_140 = 4'h8 == keyEndAddr ? io_keys_8_3_0 : _GEN_124; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_141 = 4'h8 == keyEndAddr ? io_keys_8_3_1 : _GEN_125; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_142 = 4'h8 == keyEndAddr ? io_keys_8_3_2 : _GEN_126; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_143 = 4'h8 == keyEndAddr ? io_keys_8_3_3 : _GEN_127; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_144 = 4'h9 == keyEndAddr ? io_keys_9_0_0 : _GEN_128; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_145 = 4'h9 == keyEndAddr ? io_keys_9_0_1 : _GEN_129; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_146 = 4'h9 == keyEndAddr ? io_keys_9_0_2 : _GEN_130; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_147 = 4'h9 == keyEndAddr ? io_keys_9_0_3 : _GEN_131; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_148 = 4'h9 == keyEndAddr ? io_keys_9_1_0 : _GEN_132; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_149 = 4'h9 == keyEndAddr ? io_keys_9_1_1 : _GEN_133; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_150 = 4'h9 == keyEndAddr ? io_keys_9_1_2 : _GEN_134; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_151 = 4'h9 == keyEndAddr ? io_keys_9_1_3 : _GEN_135; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_152 = 4'h9 == keyEndAddr ? io_keys_9_2_0 : _GEN_136; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_153 = 4'h9 == keyEndAddr ? io_keys_9_2_1 : _GEN_137; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_154 = 4'h9 == keyEndAddr ? io_keys_9_2_2 : _GEN_138; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_155 = 4'h9 == keyEndAddr ? io_keys_9_2_3 : _GEN_139; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_156 = 4'h9 == keyEndAddr ? io_keys_9_3_0 : _GEN_140; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_157 = 4'h9 == keyEndAddr ? io_keys_9_3_1 : _GEN_141; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_158 = 4'h9 == keyEndAddr ? io_keys_9_3_2 : _GEN_142; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_159 = 4'h9 == keyEndAddr ? io_keys_9_3_3 : _GEN_143; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_160 = 4'ha == keyEndAddr ? io_keys_10_0_0 : _GEN_144; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_161 = 4'ha == keyEndAddr ? io_keys_10_0_1 : _GEN_145; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_162 = 4'ha == keyEndAddr ? io_keys_10_0_2 : _GEN_146; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_163 = 4'ha == keyEndAddr ? io_keys_10_0_3 : _GEN_147; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_164 = 4'ha == keyEndAddr ? io_keys_10_1_0 : _GEN_148; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_165 = 4'ha == keyEndAddr ? io_keys_10_1_1 : _GEN_149; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_166 = 4'ha == keyEndAddr ? io_keys_10_1_2 : _GEN_150; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_167 = 4'ha == keyEndAddr ? io_keys_10_1_3 : _GEN_151; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_168 = 4'ha == keyEndAddr ? io_keys_10_2_0 : _GEN_152; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_169 = 4'ha == keyEndAddr ? io_keys_10_2_1 : _GEN_153; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_170 = 4'ha == keyEndAddr ? io_keys_10_2_2 : _GEN_154; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_171 = 4'ha == keyEndAddr ? io_keys_10_2_3 : _GEN_155; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_172 = 4'ha == keyEndAddr ? io_keys_10_3_0 : _GEN_156; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_173 = 4'ha == keyEndAddr ? io_keys_10_3_1 : _GEN_157; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_174 = 4'ha == keyEndAddr ? io_keys_10_3_2 : _GEN_158; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_175 = 4'ha == keyEndAddr ? io_keys_10_3_3 : _GEN_159; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_176 = 4'hb == keyEndAddr ? io_keys_11_0_0 : _GEN_160; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_177 = 4'hb == keyEndAddr ? io_keys_11_0_1 : _GEN_161; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_178 = 4'hb == keyEndAddr ? io_keys_11_0_2 : _GEN_162; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_179 = 4'hb == keyEndAddr ? io_keys_11_0_3 : _GEN_163; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_180 = 4'hb == keyEndAddr ? io_keys_11_1_0 : _GEN_164; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_181 = 4'hb == keyEndAddr ? io_keys_11_1_1 : _GEN_165; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_182 = 4'hb == keyEndAddr ? io_keys_11_1_2 : _GEN_166; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_183 = 4'hb == keyEndAddr ? io_keys_11_1_3 : _GEN_167; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_184 = 4'hb == keyEndAddr ? io_keys_11_2_0 : _GEN_168; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_185 = 4'hb == keyEndAddr ? io_keys_11_2_1 : _GEN_169; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_186 = 4'hb == keyEndAddr ? io_keys_11_2_2 : _GEN_170; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_187 = 4'hb == keyEndAddr ? io_keys_11_2_3 : _GEN_171; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_188 = 4'hb == keyEndAddr ? io_keys_11_3_0 : _GEN_172; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_189 = 4'hb == keyEndAddr ? io_keys_11_3_1 : _GEN_173; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_190 = 4'hb == keyEndAddr ? io_keys_11_3_2 : _GEN_174; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_191 = 4'hb == keyEndAddr ? io_keys_11_3_3 : _GEN_175; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_192 = 4'hc == keyEndAddr ? io_keys_12_0_0 : _GEN_176; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_193 = 4'hc == keyEndAddr ? io_keys_12_0_1 : _GEN_177; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_194 = 4'hc == keyEndAddr ? io_keys_12_0_2 : _GEN_178; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_195 = 4'hc == keyEndAddr ? io_keys_12_0_3 : _GEN_179; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_196 = 4'hc == keyEndAddr ? io_keys_12_1_0 : _GEN_180; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_197 = 4'hc == keyEndAddr ? io_keys_12_1_1 : _GEN_181; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_198 = 4'hc == keyEndAddr ? io_keys_12_1_2 : _GEN_182; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_199 = 4'hc == keyEndAddr ? io_keys_12_1_3 : _GEN_183; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_200 = 4'hc == keyEndAddr ? io_keys_12_2_0 : _GEN_184; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_201 = 4'hc == keyEndAddr ? io_keys_12_2_1 : _GEN_185; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_202 = 4'hc == keyEndAddr ? io_keys_12_2_2 : _GEN_186; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_203 = 4'hc == keyEndAddr ? io_keys_12_2_3 : _GEN_187; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_204 = 4'hc == keyEndAddr ? io_keys_12_3_0 : _GEN_188; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_205 = 4'hc == keyEndAddr ? io_keys_12_3_1 : _GEN_189; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_206 = 4'hc == keyEndAddr ? io_keys_12_3_2 : _GEN_190; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_207 = 4'hc == keyEndAddr ? io_keys_12_3_3 : _GEN_191; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_208 = 4'hd == keyEndAddr ? io_keys_13_0_0 : _GEN_192; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_209 = 4'hd == keyEndAddr ? io_keys_13_0_1 : _GEN_193; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_210 = 4'hd == keyEndAddr ? io_keys_13_0_2 : _GEN_194; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_211 = 4'hd == keyEndAddr ? io_keys_13_0_3 : _GEN_195; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_212 = 4'hd == keyEndAddr ? io_keys_13_1_0 : _GEN_196; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_213 = 4'hd == keyEndAddr ? io_keys_13_1_1 : _GEN_197; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_214 = 4'hd == keyEndAddr ? io_keys_13_1_2 : _GEN_198; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_215 = 4'hd == keyEndAddr ? io_keys_13_1_3 : _GEN_199; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_216 = 4'hd == keyEndAddr ? io_keys_13_2_0 : _GEN_200; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_217 = 4'hd == keyEndAddr ? io_keys_13_2_1 : _GEN_201; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_218 = 4'hd == keyEndAddr ? io_keys_13_2_2 : _GEN_202; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_219 = 4'hd == keyEndAddr ? io_keys_13_2_3 : _GEN_203; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_220 = 4'hd == keyEndAddr ? io_keys_13_3_0 : _GEN_204; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_221 = 4'hd == keyEndAddr ? io_keys_13_3_1 : _GEN_205; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_222 = 4'hd == keyEndAddr ? io_keys_13_3_2 : _GEN_206; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_223 = 4'hd == keyEndAddr ? io_keys_13_3_3 : _GEN_207; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_224 = 4'he == keyEndAddr ? io_keys_14_0_0 : _GEN_208; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_225 = 4'he == keyEndAddr ? io_keys_14_0_1 : _GEN_209; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_226 = 4'he == keyEndAddr ? io_keys_14_0_2 : _GEN_210; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_227 = 4'he == keyEndAddr ? io_keys_14_0_3 : _GEN_211; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_228 = 4'he == keyEndAddr ? io_keys_14_1_0 : _GEN_212; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_229 = 4'he == keyEndAddr ? io_keys_14_1_1 : _GEN_213; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_230 = 4'he == keyEndAddr ? io_keys_14_1_2 : _GEN_214; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_231 = 4'he == keyEndAddr ? io_keys_14_1_3 : _GEN_215; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_232 = 4'he == keyEndAddr ? io_keys_14_2_0 : _GEN_216; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_233 = 4'he == keyEndAddr ? io_keys_14_2_1 : _GEN_217; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_234 = 4'he == keyEndAddr ? io_keys_14_2_2 : _GEN_218; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_235 = 4'he == keyEndAddr ? io_keys_14_2_3 : _GEN_219; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_236 = 4'he == keyEndAddr ? io_keys_14_3_0 : _GEN_220; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_237 = 4'he == keyEndAddr ? io_keys_14_3_1 : _GEN_221; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_238 = 4'he == keyEndAddr ? io_keys_14_3_2 : _GEN_222; // @[AesComponents.scala 57:30]
  wire [7:0] _GEN_239 = 4'he == keyEndAddr ? io_keys_14_3_3 : _GEN_223; // @[AesComponents.scala 57:30]
  wire [7:0] xorOut_0_0 = matrix_0_0 ^ _GEN_224; // @[AesComponents.scala 57:30]
  wire [7:0] xorOut_0_1 = matrix_0_1 ^ _GEN_225; // @[AesComponents.scala 57:51]
  wire [7:0] xorOut_0_2 = matrix_0_2 ^ _GEN_226; // @[AesComponents.scala 57:72]
  wire [7:0] xorOut_0_3 = matrix_0_3 ^ _GEN_227; // @[AesComponents.scala 57:93]
  wire [7:0] xorOut_1_0 = matrix_1_0 ^ _GEN_228; // @[AesComponents.scala 58:30]
  wire [7:0] xorOut_1_1 = matrix_1_1 ^ _GEN_229; // @[AesComponents.scala 58:51]
  wire [7:0] xorOut_1_2 = matrix_1_2 ^ _GEN_230; // @[AesComponents.scala 58:72]
  wire [7:0] xorOut_1_3 = matrix_1_3 ^ _GEN_231; // @[AesComponents.scala 58:93]
  wire [7:0] xorOut_2_0 = matrix_2_0 ^ _GEN_232; // @[AesComponents.scala 59:30]
  wire [7:0] xorOut_2_1 = matrix_2_1 ^ _GEN_233; // @[AesComponents.scala 59:51]
  wire [7:0] xorOut_2_2 = matrix_2_2 ^ _GEN_234; // @[AesComponents.scala 59:72]
  wire [7:0] xorOut_2_3 = matrix_2_3 ^ _GEN_235; // @[AesComponents.scala 59:93]
  wire [7:0] xorOut_3_0 = matrix_3_0 ^ _GEN_236; // @[AesComponents.scala 60:30]
  wire [7:0] xorOut_3_1 = matrix_3_1 ^ _GEN_237; // @[AesComponents.scala 60:51]
  wire [7:0] xorOut_3_2 = matrix_3_2 ^ _GEN_238; // @[AesComponents.scala 60:72]
  wire [7:0] xorOut_3_3 = matrix_3_3 ^ _GEN_239; // @[AesComponents.scala 60:93]
  wire [7:0] _T_4534 = xorOut_0_0 ^ xorOut_0_2; // @[AesComponents.scala 100:47]
  wire [7:0] _T_4535 = _T_4534 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4536 = _T_4535 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4537 = {_T_4534, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4538 = _T_4537 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4539 = _T_4538 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4541 = _T_4536 ? _T_4539 : _T_4537; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4542 = _T_4541 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4543 = _T_4542 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4544 = {_T_4541, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4545 = _T_4544 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4546 = _T_4545 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4548 = _T_4543 ? _T_4546 : _T_4544; // @[AesComponents.scala 88:38]
  wire [7:0] _T_4549 = xorOut_0_1 ^ xorOut_0_3; // @[AesComponents.scala 101:47]
  wire [7:0] _T_4550 = _T_4549 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4551 = _T_4550 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4552 = {_T_4549, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4553 = _T_4552 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4554 = _T_4553 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4556 = _T_4551 ? _T_4554 : _T_4552; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4557 = _T_4556 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4558 = _T_4557 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4559 = {_T_4556, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4560 = _T_4559 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4561 = _T_4560 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4563 = _T_4558 ? _T_4561 : _T_4559; // @[AesComponents.scala 88:38]
  wire [9:0] _GEN_311 = {{2'd0}, xorOut_0_0}; // @[AesComponents.scala 102:34]
  wire [9:0] _T_4564 = _GEN_311 ^ _T_4548; // @[AesComponents.scala 102:34]
  wire [9:0] _GEN_312 = {{2'd0}, xorOut_0_1}; // @[AesComponents.scala 103:34]
  wire [9:0] _T_4565 = _GEN_312 ^ _T_4563; // @[AesComponents.scala 103:34]
  wire [9:0] _GEN_313 = {{2'd0}, xorOut_0_2}; // @[AesComponents.scala 104:34]
  wire [9:0] _T_4566 = _GEN_313 ^ _T_4548; // @[AesComponents.scala 104:34]
  wire [9:0] _GEN_314 = {{2'd0}, xorOut_0_3}; // @[AesComponents.scala 105:34]
  wire [9:0] _T_4567 = _GEN_314 ^ _T_4563; // @[AesComponents.scala 105:34]
  wire [7:0] _T_4568 = xorOut_1_0 ^ xorOut_1_2; // @[AesComponents.scala 100:47]
  wire [7:0] _T_4569 = _T_4568 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4570 = _T_4569 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4571 = {_T_4568, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4572 = _T_4571 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4573 = _T_4572 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4575 = _T_4570 ? _T_4573 : _T_4571; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4576 = _T_4575 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4577 = _T_4576 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4578 = {_T_4575, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4579 = _T_4578 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4580 = _T_4579 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4582 = _T_4577 ? _T_4580 : _T_4578; // @[AesComponents.scala 88:38]
  wire [7:0] _T_4583 = xorOut_1_1 ^ xorOut_1_3; // @[AesComponents.scala 101:47]
  wire [7:0] _T_4584 = _T_4583 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4585 = _T_4584 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4586 = {_T_4583, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4587 = _T_4586 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4588 = _T_4587 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4590 = _T_4585 ? _T_4588 : _T_4586; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4591 = _T_4590 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4592 = _T_4591 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4593 = {_T_4590, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4594 = _T_4593 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4595 = _T_4594 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4597 = _T_4592 ? _T_4595 : _T_4593; // @[AesComponents.scala 88:38]
  wire [9:0] _GEN_315 = {{2'd0}, xorOut_1_0}; // @[AesComponents.scala 102:34]
  wire [9:0] _T_4598 = _GEN_315 ^ _T_4582; // @[AesComponents.scala 102:34]
  wire [9:0] _GEN_316 = {{2'd0}, xorOut_1_1}; // @[AesComponents.scala 103:34]
  wire [9:0] _T_4599 = _GEN_316 ^ _T_4597; // @[AesComponents.scala 103:34]
  wire [9:0] _GEN_317 = {{2'd0}, xorOut_1_2}; // @[AesComponents.scala 104:34]
  wire [9:0] _T_4600 = _GEN_317 ^ _T_4582; // @[AesComponents.scala 104:34]
  wire [9:0] _GEN_318 = {{2'd0}, xorOut_1_3}; // @[AesComponents.scala 105:34]
  wire [9:0] _T_4601 = _GEN_318 ^ _T_4597; // @[AesComponents.scala 105:34]
  wire [7:0] _T_4602 = xorOut_2_0 ^ xorOut_2_2; // @[AesComponents.scala 100:47]
  wire [7:0] _T_4603 = _T_4602 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4604 = _T_4603 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4605 = {_T_4602, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4606 = _T_4605 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4607 = _T_4606 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4609 = _T_4604 ? _T_4607 : _T_4605; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4610 = _T_4609 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4611 = _T_4610 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4612 = {_T_4609, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4613 = _T_4612 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4614 = _T_4613 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4616 = _T_4611 ? _T_4614 : _T_4612; // @[AesComponents.scala 88:38]
  wire [7:0] _T_4617 = xorOut_2_1 ^ xorOut_2_3; // @[AesComponents.scala 101:47]
  wire [7:0] _T_4618 = _T_4617 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4619 = _T_4618 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4620 = {_T_4617, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4621 = _T_4620 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4622 = _T_4621 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4624 = _T_4619 ? _T_4622 : _T_4620; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4625 = _T_4624 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4626 = _T_4625 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4627 = {_T_4624, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4628 = _T_4627 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4629 = _T_4628 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4631 = _T_4626 ? _T_4629 : _T_4627; // @[AesComponents.scala 88:38]
  wire [9:0] _GEN_319 = {{2'd0}, xorOut_2_0}; // @[AesComponents.scala 102:34]
  wire [9:0] _T_4632 = _GEN_319 ^ _T_4616; // @[AesComponents.scala 102:34]
  wire [9:0] _GEN_320 = {{2'd0}, xorOut_2_1}; // @[AesComponents.scala 103:34]
  wire [9:0] _T_4633 = _GEN_320 ^ _T_4631; // @[AesComponents.scala 103:34]
  wire [9:0] _GEN_321 = {{2'd0}, xorOut_2_2}; // @[AesComponents.scala 104:34]
  wire [9:0] _T_4634 = _GEN_321 ^ _T_4616; // @[AesComponents.scala 104:34]
  wire [9:0] _GEN_322 = {{2'd0}, xorOut_2_3}; // @[AesComponents.scala 105:34]
  wire [9:0] _T_4635 = _GEN_322 ^ _T_4631; // @[AesComponents.scala 105:34]
  wire [7:0] _T_4636 = xorOut_3_0 ^ xorOut_3_2; // @[AesComponents.scala 100:47]
  wire [7:0] _T_4637 = _T_4636 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4638 = _T_4637 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4639 = {_T_4636, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4640 = _T_4639 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4641 = _T_4640 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4643 = _T_4638 ? _T_4641 : _T_4639; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4644 = _T_4643 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4645 = _T_4644 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4646 = {_T_4643, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4647 = _T_4646 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4648 = _T_4647 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4650 = _T_4645 ? _T_4648 : _T_4646; // @[AesComponents.scala 88:38]
  wire [7:0] _T_4651 = xorOut_3_1 ^ xorOut_3_3; // @[AesComponents.scala 101:47]
  wire [7:0] _T_4652 = _T_4651 & 8'h80; // @[AesComponents.scala 88:42]
  wire  _T_4653 = _T_4652 != 8'h0; // @[AesComponents.scala 88:52]
  wire [8:0] _T_4654 = {_T_4651, 1'h0}; // @[AesComponents.scala 88:65]
  wire [8:0] _T_4655 = _T_4654 ^ 9'h1b; // @[AesComponents.scala 88:78]
  wire [8:0] _T_4656 = _T_4655 & 9'hff; // @[AesComponents.scala 88:88]
  wire [8:0] _T_4658 = _T_4653 ? _T_4656 : _T_4654; // @[AesComponents.scala 88:38]
  wire [8:0] _T_4659 = _T_4658 & 9'h80; // @[AesComponents.scala 88:42]
  wire  _T_4660 = _T_4659 != 9'h0; // @[AesComponents.scala 88:52]
  wire [9:0] _T_4661 = {_T_4658, 1'h0}; // @[AesComponents.scala 88:65]
  wire [9:0] _T_4662 = _T_4661 ^ 10'h1b; // @[AesComponents.scala 88:78]
  wire [9:0] _T_4663 = _T_4662 & 10'hff; // @[AesComponents.scala 88:88]
  wire [9:0] _T_4665 = _T_4660 ? _T_4663 : _T_4661; // @[AesComponents.scala 88:38]
  wire [9:0] _GEN_323 = {{2'd0}, xorOut_3_0}; // @[AesComponents.scala 102:34]
  wire [9:0] _T_4666 = _GEN_323 ^ _T_4650; // @[AesComponents.scala 102:34]
  wire [9:0] _GEN_324 = {{2'd0}, xorOut_3_1}; // @[AesComponents.scala 103:34]
  wire [9:0] _T_4667 = _GEN_324 ^ _T_4665; // @[AesComponents.scala 103:34]
  wire [9:0] _GEN_325 = {{2'd0}, xorOut_3_2}; // @[AesComponents.scala 104:34]
  wire [9:0] _T_4668 = _GEN_325 ^ _T_4650; // @[AesComponents.scala 104:34]
  wire [9:0] _GEN_326 = {{2'd0}, xorOut_3_3}; // @[AesComponents.scala 105:34]
  wire [9:0] _T_4669 = _GEN_326 ^ _T_4665; // @[AesComponents.scala 105:34]
  wire [63:0] _T_4717 = {xorOut_2_0,xorOut_2_1,xorOut_2_2,xorOut_2_3,xorOut_3_0,xorOut_3_1,xorOut_3_2,xorOut_3_3}; // @[Cat.scala 29:58]
  wire [127:0] _T_4725 = {xorOut_0_0,xorOut_0_1,xorOut_0_2,xorOut_0_3,xorOut_1_0,xorOut_1_1,xorOut_1_2,xorOut_1_3,_T_4717}; // @[Cat.scala 29:58]
  wire [127:0] _T_4726 = io_ivIn ^ _T_4725; // @[AesDecrypt.scala 79:37]
  wire [7:0] finalOut_0_0 = _T_4726[127:120]; // @[AesComponents.scala 43:25]
  wire [7:0] finalOut_0_1 = _T_4726[119:112]; // @[AesComponents.scala 43:45]
  wire [7:0] finalOut_0_2 = _T_4726[111:104]; // @[AesComponents.scala 43:65]
  wire [7:0] finalOut_0_3 = _T_4726[103:96]; // @[AesComponents.scala 43:85]
  wire [7:0] finalOut_1_0 = _T_4726[95:88]; // @[AesComponents.scala 44:25]
  wire [7:0] finalOut_1_1 = _T_4726[87:80]; // @[AesComponents.scala 44:45]
  wire [7:0] finalOut_1_2 = _T_4726[79:72]; // @[AesComponents.scala 44:65]
  wire [7:0] finalOut_1_3 = _T_4726[71:64]; // @[AesComponents.scala 44:85]
  wire [7:0] finalOut_2_0 = _T_4726[63:56]; // @[AesComponents.scala 45:25]
  wire [7:0] finalOut_2_1 = _T_4726[55:48]; // @[AesComponents.scala 45:45]
  wire [7:0] finalOut_2_2 = _T_4726[47:40]; // @[AesComponents.scala 45:65]
  wire [7:0] finalOut_2_3 = _T_4726[39:32]; // @[AesComponents.scala 45:85]
  wire [7:0] finalOut_3_0 = _T_4726[31:24]; // @[AesComponents.scala 46:25]
  wire [7:0] finalOut_3_1 = _T_4726[23:16]; // @[AesComponents.scala 46:45]
  wire [7:0] finalOut_3_2 = _T_4726[15:8]; // @[AesComponents.scala 46:65]
  wire [7:0] finalOut_3_3 = _T_4726[7:0]; // @[AesComponents.scala 46:85]
  wire  _T_4747 = io_ready & io_dataValid; // @[AesDecrypt.scala 81:20]
  wire [4:0] _T_4769 = io_aes256 ? 5'h1d : 5'h15; // @[AesDecrypt.scala 85:21]
  wire  _T_4770 = ~io_ready; // @[AesDecrypt.scala 88:11]
  wire  _T_4771 = state == 6'h1; // @[AesDecrypt.scala 89:21]
  wire  _T_4773 = ~state[0]; // @[AesDecrypt.scala 92:31]
  wire [5:0] _GEN_327 = {{1'd0}, _T_4769}; // @[AesDecrypt.scala 95:33]
  wire  _T_4775 = state == _GEN_327; // @[AesDecrypt.scala 95:33]
  wire  _GEN_275 = _T_4773 ? 1'h0 : 1'h1; // @[AesDecrypt.scala 92:40]
  wire  _GEN_292 = _T_4771 | _GEN_275; // @[AesDecrypt.scala 89:30]
  wire [5:0] _T_4778 = state - 6'h1; // @[AesDecrypt.scala 99:24]
  MixColsModule MixColsModule ( // @[AesComponents.scala 91:35]
    .io_in_0_0(MixColsModule_io_in_0_0),
    .io_in_0_1(MixColsModule_io_in_0_1),
    .io_in_0_2(MixColsModule_io_in_0_2),
    .io_in_0_3(MixColsModule_io_in_0_3),
    .io_in_1_0(MixColsModule_io_in_1_0),
    .io_in_1_1(MixColsModule_io_in_1_1),
    .io_in_1_2(MixColsModule_io_in_1_2),
    .io_in_1_3(MixColsModule_io_in_1_3),
    .io_in_2_0(MixColsModule_io_in_2_0),
    .io_in_2_1(MixColsModule_io_in_2_1),
    .io_in_2_2(MixColsModule_io_in_2_2),
    .io_in_2_3(MixColsModule_io_in_2_3),
    .io_in_3_0(MixColsModule_io_in_3_0),
    .io_in_3_1(MixColsModule_io_in_3_1),
    .io_in_3_2(MixColsModule_io_in_3_2),
    .io_in_3_3(MixColsModule_io_in_3_3),
    .io_out_0_0(MixColsModule_io_out_0_0),
    .io_out_0_1(MixColsModule_io_out_0_1),
    .io_out_0_2(MixColsModule_io_out_0_2),
    .io_out_0_3(MixColsModule_io_out_0_3),
    .io_out_1_0(MixColsModule_io_out_1_0),
    .io_out_1_1(MixColsModule_io_out_1_1),
    .io_out_1_2(MixColsModule_io_out_1_2),
    .io_out_1_3(MixColsModule_io_out_1_3),
    .io_out_2_0(MixColsModule_io_out_2_0),
    .io_out_2_1(MixColsModule_io_out_2_1),
    .io_out_2_2(MixColsModule_io_out_2_2),
    .io_out_2_3(MixColsModule_io_out_2_3),
    .io_out_3_0(MixColsModule_io_out_3_0),
    .io_out_3_1(MixColsModule_io_out_3_1),
    .io_out_3_2(MixColsModule_io_out_3_2),
    .io_out_3_3(MixColsModule_io_out_3_3)
  );
  assign io_shiftCyc = io_shift; // @[AesDecrypt.scala 59:17]
  assign io_shiftRev = io_shift; // @[AesDecrypt.scala 58:17]
  assign io_shift = _T_4770 & _GEN_292; // @[AesDecrypt.scala 60:14 AesDecrypt.scala 91:22 AesDecrypt.scala 96:22]
  assign io_ready = _T | _T_1; // @[AesDecrypt.scala 55:14]
  assign io_dataOut = {_T_17,_T_10}; // @[AesDecrypt.scala 67:16]
  assign io_ivOut = ctSaved; // @[AesDecrypt.scala 68:14]
  assign io_outputValid = state == 6'h0; // @[AesDecrypt.scala 56:20]
  assign MixColsModule_io_in_0_0 = _T_4564[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_0_1 = _T_4565[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_0_2 = _T_4566[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_0_3 = _T_4567[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_0 = _T_4598[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_1 = _T_4599[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_2 = _T_4600[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_1_3 = _T_4601[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_0 = _T_4632[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_1 = _T_4633[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_2 = _T_4634[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_2_3 = _T_4635[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_0 = _T_4666[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_1 = _T_4667[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_2 = _T_4668[7:0]; // @[AesComponents.scala 92:29]
  assign MixColsModule_io_in_3_3 = _T_4669[7:0]; // @[AesComponents.scala 92:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[5:0];
  _RAND_1 = {4{`RANDOM}};
  ctSaved = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  matrix_0_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  matrix_0_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  matrix_0_2 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  matrix_0_3 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  matrix_1_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  matrix_1_1 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  matrix_1_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  matrix_1_3 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  matrix_2_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  matrix_2_1 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  matrix_2_2 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  matrix_2_3 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  matrix_3_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  matrix_3_1 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  matrix_3_2 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  matrix_3_3 = _RAND_17[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 6'h1e;
    end else if (_T_4770) begin
      state <= _T_4778;
    end else if (_T_4747) begin
      state <= {{1'd0}, _T_4769};
    end
    if (_T_4747) begin
      ctSaved <= io_dataIn;
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_0_0 <= finalOut_0_0;
      end else if (_T_4773) begin
        matrix_0_0 <= roundPart1_0_0;
      end else if (_T_4775) begin
        matrix_0_0 <= xorOut_0_0;
      end else begin
        matrix_0_0 <= MixColsModule_io_out_0_0;
      end
    end else if (_T_4747) begin
      matrix_0_0 <= io_dataIn[127:120];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_0_1 <= finalOut_0_1;
      end else if (_T_4773) begin
        matrix_0_1 <= roundPart1_0_1;
      end else if (_T_4775) begin
        matrix_0_1 <= xorOut_0_1;
      end else begin
        matrix_0_1 <= MixColsModule_io_out_0_1;
      end
    end else if (_T_4747) begin
      matrix_0_1 <= io_dataIn[119:112];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_0_2 <= finalOut_0_2;
      end else if (_T_4773) begin
        matrix_0_2 <= roundPart1_0_2;
      end else if (_T_4775) begin
        matrix_0_2 <= xorOut_0_2;
      end else begin
        matrix_0_2 <= MixColsModule_io_out_0_2;
      end
    end else if (_T_4747) begin
      matrix_0_2 <= io_dataIn[111:104];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_0_3 <= finalOut_0_3;
      end else if (_T_4773) begin
        matrix_0_3 <= roundPart1_0_3;
      end else if (_T_4775) begin
        matrix_0_3 <= xorOut_0_3;
      end else begin
        matrix_0_3 <= MixColsModule_io_out_0_3;
      end
    end else if (_T_4747) begin
      matrix_0_3 <= io_dataIn[103:96];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_1_0 <= finalOut_1_0;
      end else if (_T_4773) begin
        matrix_1_0 <= roundPart1_1_0;
      end else if (_T_4775) begin
        matrix_1_0 <= xorOut_1_0;
      end else begin
        matrix_1_0 <= MixColsModule_io_out_1_0;
      end
    end else if (_T_4747) begin
      matrix_1_0 <= io_dataIn[95:88];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_1_1 <= finalOut_1_1;
      end else if (_T_4773) begin
        matrix_1_1 <= roundPart1_1_1;
      end else if (_T_4775) begin
        matrix_1_1 <= xorOut_1_1;
      end else begin
        matrix_1_1 <= MixColsModule_io_out_1_1;
      end
    end else if (_T_4747) begin
      matrix_1_1 <= io_dataIn[87:80];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_1_2 <= finalOut_1_2;
      end else if (_T_4773) begin
        matrix_1_2 <= roundPart1_1_2;
      end else if (_T_4775) begin
        matrix_1_2 <= xorOut_1_2;
      end else begin
        matrix_1_2 <= MixColsModule_io_out_1_2;
      end
    end else if (_T_4747) begin
      matrix_1_2 <= io_dataIn[79:72];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_1_3 <= finalOut_1_3;
      end else if (_T_4773) begin
        matrix_1_3 <= roundPart1_1_3;
      end else if (_T_4775) begin
        matrix_1_3 <= xorOut_1_3;
      end else begin
        matrix_1_3 <= MixColsModule_io_out_1_3;
      end
    end else if (_T_4747) begin
      matrix_1_3 <= io_dataIn[71:64];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_2_0 <= finalOut_2_0;
      end else if (_T_4773) begin
        matrix_2_0 <= roundPart1_2_0;
      end else if (_T_4775) begin
        matrix_2_0 <= xorOut_2_0;
      end else begin
        matrix_2_0 <= MixColsModule_io_out_2_0;
      end
    end else if (_T_4747) begin
      matrix_2_0 <= io_dataIn[63:56];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_2_1 <= finalOut_2_1;
      end else if (_T_4773) begin
        matrix_2_1 <= roundPart1_2_1;
      end else if (_T_4775) begin
        matrix_2_1 <= xorOut_2_1;
      end else begin
        matrix_2_1 <= MixColsModule_io_out_2_1;
      end
    end else if (_T_4747) begin
      matrix_2_1 <= io_dataIn[55:48];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_2_2 <= finalOut_2_2;
      end else if (_T_4773) begin
        matrix_2_2 <= roundPart1_2_2;
      end else if (_T_4775) begin
        matrix_2_2 <= xorOut_2_2;
      end else begin
        matrix_2_2 <= MixColsModule_io_out_2_2;
      end
    end else if (_T_4747) begin
      matrix_2_2 <= io_dataIn[47:40];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_2_3 <= finalOut_2_3;
      end else if (_T_4773) begin
        matrix_2_3 <= roundPart1_2_3;
      end else if (_T_4775) begin
        matrix_2_3 <= xorOut_2_3;
      end else begin
        matrix_2_3 <= MixColsModule_io_out_2_3;
      end
    end else if (_T_4747) begin
      matrix_2_3 <= io_dataIn[39:32];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_3_0 <= finalOut_3_0;
      end else if (_T_4773) begin
        matrix_3_0 <= roundPart1_3_0;
      end else if (_T_4775) begin
        matrix_3_0 <= xorOut_3_0;
      end else begin
        matrix_3_0 <= MixColsModule_io_out_3_0;
      end
    end else if (_T_4747) begin
      matrix_3_0 <= io_dataIn[31:24];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_3_1 <= finalOut_3_1;
      end else if (_T_4773) begin
        matrix_3_1 <= roundPart1_3_1;
      end else if (_T_4775) begin
        matrix_3_1 <= xorOut_3_1;
      end else begin
        matrix_3_1 <= MixColsModule_io_out_3_1;
      end
    end else if (_T_4747) begin
      matrix_3_1 <= io_dataIn[23:16];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_3_2 <= finalOut_3_2;
      end else if (_T_4773) begin
        matrix_3_2 <= roundPart1_3_2;
      end else if (_T_4775) begin
        matrix_3_2 <= xorOut_3_2;
      end else begin
        matrix_3_2 <= MixColsModule_io_out_3_2;
      end
    end else if (_T_4747) begin
      matrix_3_2 <= io_dataIn[15:8];
    end
    if (_T_4770) begin
      if (_T_4771) begin
        matrix_3_3 <= finalOut_3_3;
      end else if (_T_4773) begin
        matrix_3_3 <= roundPart1_3_3;
      end else if (_T_4775) begin
        matrix_3_3 <= xorOut_3_3;
      end else begin
        matrix_3_3 <= MixColsModule_io_out_3_3;
      end
    end else if (_T_4747) begin
      matrix_3_3 <= io_dataIn[7:0];
    end
  end
endmodule
module AesCombined(
  input          clock,
  input          reset,
  input  [127:0] io_encDataIn,
  input  [127:0] io_encIvIn,
  input          io_encDataValid,
  input  [127:0] io_decDataIn,
  input  [127:0] io_decIvIn,
  input          io_decDataValid,
  input          io_aes256,
  input  [127:0] io_keyIn,
  input          io_keyShift,
  input          io_keyValid,
  output         io_encReady,
  output         io_decReady,
  output [127:0] io_encDataOut,
  output [127:0] io_encIvOut,
  output         io_encOutputValid,
  output [127:0] io_decDataOut,
  output [127:0] io_decIvOut,
  output         io_decOutputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  shreg_clock; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_input; // @[AesCombined.scala 55:23]
  wire  shreg_io_enable; // @[AesCombined.scala 55:23]
  wire  shreg_io_rev; // @[AesCombined.scala 55:23]
  wire  shreg_io_cyc; // @[AesCombined.scala 55:23]
  wire  shreg_io_tap; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_0; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_1; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_2; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_3; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_4; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_5; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_6; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_7; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_8; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_9; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_10; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_11; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_12; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_13; // @[AesCombined.scala 55:23]
  wire [127:0] shreg_io_output_14; // @[AesCombined.scala 55:23]
  wire  enc_clock; // @[AesCombined.scala 84:21]
  wire  enc_reset; // @[AesCombined.scala 84:21]
  wire [127:0] enc_io_dataIn; // @[AesCombined.scala 84:21]
  wire [127:0] enc_io_ivIn; // @[AesCombined.scala 84:21]
  wire  enc_io_dataValid; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_0_0; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_0_1; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_0_2; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_0_3; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_1_0; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_1_1; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_1_2; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_1_3; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_2_0; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_2_1; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_2_2; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_2_3; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_3_0; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_3_1; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_3_2; // @[AesCombined.scala 84:21]
  wire [7:0] enc_io_keys_0_3_3; // @[AesCombined.scala 84:21]
  wire  enc_io_aes256; // @[AesCombined.scala 84:21]
  wire  enc_io_shiftCyc; // @[AesCombined.scala 84:21]
  wire  enc_io_shift; // @[AesCombined.scala 84:21]
  wire  enc_io_ready; // @[AesCombined.scala 84:21]
  wire [127:0] enc_io_dataOut; // @[AesCombined.scala 84:21]
  wire [127:0] enc_io_ivOut; // @[AesCombined.scala 84:21]
  wire  enc_io_outputValid; // @[AesCombined.scala 84:21]
  wire  dec_clock; // @[AesCombined.scala 97:21]
  wire  dec_reset; // @[AesCombined.scala 97:21]
  wire [127:0] dec_io_dataIn; // @[AesCombined.scala 97:21]
  wire [127:0] dec_io_ivIn; // @[AesCombined.scala 97:21]
  wire  dec_io_dataValid; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_0_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_1_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_2_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_3_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_4_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_5_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_6_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_7_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_8_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_9_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_10_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_11_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_12_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_13_3_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_0_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_0_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_0_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_0_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_1_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_1_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_1_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_1_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_2_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_2_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_2_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_2_3; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_3_0; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_3_1; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_3_2; // @[AesCombined.scala 97:21]
  wire [7:0] dec_io_keys_14_3_3; // @[AesCombined.scala 97:21]
  wire  dec_io_aes256; // @[AesCombined.scala 97:21]
  wire  dec_io_shiftCyc; // @[AesCombined.scala 97:21]
  wire  dec_io_shiftRev; // @[AesCombined.scala 97:21]
  wire  dec_io_shift; // @[AesCombined.scala 97:21]
  wire  dec_io_ready; // @[AesCombined.scala 97:21]
  wire [127:0] dec_io_dataOut; // @[AesCombined.scala 97:21]
  wire [127:0] dec_io_ivOut; // @[AesCombined.scala 97:21]
  wire  dec_io_outputValid; // @[AesCombined.scala 97:21]
  reg  keyUpdate; // @[AesCombined.scala 52:28]
  reg [5:0] keyInd; // @[AesCombined.scala 53:25]
  wire  _GEN_0 = io_keyValid | keyUpdate; // @[AesCombined.scala 61:24]
  wire  _T = io_keyValid | io_keyShift; // @[AesCombined.scala 66:23]
  wire [127:0] _GEN_3 = _T ? io_keyIn : 128'h0; // @[AesCombined.scala 66:39]
  wire [5:0] _T_2 = keyInd + 6'h1; // @[AesCombined.scala 72:26]
  wire [3:0] _T_5 = io_aes256 ? 4'he : 4'hf; // @[AesCombined.scala 74:35]
  wire [5:0] _GEN_42 = {{2'd0}, _T_5}; // @[AesCombined.scala 74:28]
  wire  _T_6 = _T_2 == _GEN_42; // @[AesCombined.scala 74:28]
  wire  _T_51 = ~keyInd[0]; // @[AesComponents.scala 114:25]
  wire  _T_52 = _T_51 & io_aes256; // @[AesComponents.scala 114:38]
  wire  _T_70 = shreg_io_output_0[25] ^ shreg_io_output_0[27]; // @[AesSbox.scala 40:63]
  wire  _T_72 = shreg_io_output_0[28] ^ shreg_io_output_0[31]; // @[AesSbox.scala 40:63]
  wire  _T_74 = shreg_io_output_0[30] ^ shreg_io_output_0[29]; // @[AesSbox.scala 40:63]
  wire  _T_76 = shreg_io_output_0[24] ^ _T_74; // @[AesSbox.scala 40:63]
  wire  _T_78 = _T_70 ^ _T_72; // @[AesSbox.scala 40:63]
  wire  _T_80 = shreg_io_output_0[30] ^ shreg_io_output_0[26]; // @[AesSbox.scala 40:63]
  wire  _T_82 = shreg_io_output_0[31] ^ shreg_io_output_0[25]; // @[AesSbox.scala 40:63]
  wire  _T_84 = _T_70 ^ _T_80; // @[AesSbox.scala 40:63]
  wire  _T_86 = shreg_io_output_0[25] ^ _T_76; // @[AesSbox.scala 40:63]
  wire  _T_88 = shreg_io_output_0[28] ^ _T_76; // @[AesSbox.scala 40:63]
  wire  _T_90 = shreg_io_output_0[24] ^ _T_78; // @[AesSbox.scala 40:63]
  wire  _T_92 = _T_78 ^ _T_80; // @[AesSbox.scala 40:63]
  wire  _T_94 = shreg_io_output_0[29] ^ shreg_io_output_0[26]; // @[AesSbox.scala 40:63]
  wire  _T_96 = _T_74 ^ _T_78; // @[AesSbox.scala 40:63]
  wire  _T_98 = shreg_io_output_0[26] ^ _T_82; // @[AesSbox.scala 40:63]
  wire  _T_100 = shreg_io_output_0[31] ^ shreg_io_output_0[26]; // @[AesSbox.scala 40:63]
  wire  _T_102 = shreg_io_output_0[24] ^ _T_84; // @[AesSbox.scala 40:63]
  wire  _T_104 = shreg_io_output_0[25] ^ shreg_io_output_0[26]; // @[AesSbox.scala 40:63]
  wire  _T_106 = _T_72 ^ _T_104; // @[AesSbox.scala 40:63]
  wire  _T_108 = _T_76 ^ _T_98; // @[AesSbox.scala 40:63]
  wire  _T_110 = _T_70 ^ _T_94; // @[AesSbox.scala 40:63]
  wire  _T_112 = shreg_io_output_0[31] ^ _T_76; // @[AesSbox.scala 40:63]
  wire  _T_114 = _T_110 ^ _T_78; // @[AesSbox.scala 40:63]
  wire  _T_116 = _T_110 ^ _T_82; // @[AesSbox.scala 40:63]
  wire  _T_118 = _T_82 ^ _T_106; // @[AesSbox.scala 40:63]
  wire  _T_120 = _T_100 ^ _T_96; // @[AesSbox.scala 40:63]
  wire  _T_122 = _T_112 ^ _T_102; // @[AesSbox.scala 40:63]
  wire  _T_124 = _T_106 & _T_78; // @[AesSbox.scala 41:63]
  wire  _T_126 = _T_108 & _T_90; // @[AesSbox.scala 41:63]
  wire  _T_128 = _T_92 ^ _T_124; // @[AesSbox.scala 40:63]
  wire  _T_130 = _T_88 & shreg_io_output_0[24]; // @[AesSbox.scala 41:63]
  wire  _T_132 = _T_130 ^ _T_124; // @[AesSbox.scala 40:63]
  wire  _T_134 = _T_82 & _T_110; // @[AesSbox.scala 41:63]
  wire  _T_136 = _T_86 & _T_76; // @[AesSbox.scala 41:63]
  wire  _T_138 = _T_116 ^ _T_134; // @[AesSbox.scala 40:63]
  wire  _T_140 = _T_112 & _T_102; // @[AesSbox.scala 41:63]
  wire  _T_142 = _T_140 ^ _T_134; // @[AesSbox.scala 40:63]
  wire  _T_144 = _T_72 & _T_84; // @[AesSbox.scala 41:63]
  wire  _T_146 = _T_118 & _T_114; // @[AesSbox.scala 41:63]
  wire  _T_148 = _T_146 ^ _T_144; // @[AesSbox.scala 40:63]
  wire  _T_150 = _T_100 & _T_96; // @[AesSbox.scala 41:63]
  wire  _T_152 = _T_150 ^ _T_144; // @[AesSbox.scala 40:63]
  wire  _T_154 = _T_128 ^ _T_126; // @[AesSbox.scala 40:63]
  wire  _T_156 = _T_132 ^ _T_120; // @[AesSbox.scala 40:63]
  wire  _T_158 = _T_138 ^ _T_136; // @[AesSbox.scala 40:63]
  wire  _T_160 = _T_142 ^ _T_152; // @[AesSbox.scala 40:63]
  wire  _T_162 = _T_154 ^ _T_148; // @[AesSbox.scala 40:63]
  wire  _T_164 = _T_156 ^ _T_152; // @[AesSbox.scala 40:63]
  wire  _T_166 = _T_158 ^ _T_148; // @[AesSbox.scala 40:63]
  wire  _T_168 = _T_160 ^ _T_122; // @[AesSbox.scala 40:63]
  wire  _T_170 = _T_166 ^ _T_168; // @[AesSbox.scala 40:63]
  wire  _T_172 = _T_166 & _T_162; // @[AesSbox.scala 41:63]
  wire  _T_174 = _T_164 ^ _T_172; // @[AesSbox.scala 40:63]
  wire  _T_176 = _T_162 ^ _T_164; // @[AesSbox.scala 40:63]
  wire  _T_178 = _T_168 ^ _T_172; // @[AesSbox.scala 40:63]
  wire  _T_180 = _T_178 & _T_176; // @[AesSbox.scala 41:63]
  wire  _T_182 = _T_174 & _T_170; // @[AesSbox.scala 41:63]
  wire  _T_184 = _T_162 & _T_168; // @[AesSbox.scala 41:63]
  wire  _T_186 = _T_176 & _T_184; // @[AesSbox.scala 41:63]
  wire  _T_188 = _T_176 ^ _T_172; // @[AesSbox.scala 40:63]
  wire  _T_190 = _T_164 & _T_166; // @[AesSbox.scala 41:63]
  wire  _T_192 = _T_170 & _T_190; // @[AesSbox.scala 41:63]
  wire  _T_194 = _T_170 ^ _T_172; // @[AesSbox.scala 40:63]
  wire  _T_196 = _T_164 ^ _T_180; // @[AesSbox.scala 40:63]
  wire  _T_198 = _T_186 ^ _T_188; // @[AesSbox.scala 40:63]
  wire  _T_200 = _T_168 ^ _T_182; // @[AesSbox.scala 40:63]
  wire  _T_202 = _T_192 ^ _T_194; // @[AesSbox.scala 40:63]
  wire  _T_204 = _T_198 ^ _T_202; // @[AesSbox.scala 40:63]
  wire  _T_206 = _T_196 ^ _T_200; // @[AesSbox.scala 40:63]
  wire  _T_208 = _T_196 ^ _T_198; // @[AesSbox.scala 40:63]
  wire  _T_210 = _T_200 ^ _T_202; // @[AesSbox.scala 40:63]
  wire  _T_212 = _T_206 ^ _T_204; // @[AesSbox.scala 40:63]
  wire  _T_214 = _T_210 & _T_78; // @[AesSbox.scala 41:63]
  wire  _T_216 = _T_202 & _T_90; // @[AesSbox.scala 41:63]
  wire  _T_218 = _T_200 & shreg_io_output_0[24]; // @[AesSbox.scala 41:63]
  wire  _T_220 = _T_208 & _T_110; // @[AesSbox.scala 41:63]
  wire  _T_222 = _T_198 & _T_76; // @[AesSbox.scala 41:63]
  wire  _T_224 = _T_196 & _T_102; // @[AesSbox.scala 41:63]
  wire  _T_226 = _T_206 & _T_84; // @[AesSbox.scala 41:63]
  wire  _T_228 = _T_212 & _T_114; // @[AesSbox.scala 41:63]
  wire  _T_230 = _T_204 & _T_96; // @[AesSbox.scala 41:63]
  wire  _T_232 = _T_210 & _T_106; // @[AesSbox.scala 41:63]
  wire  _T_234 = _T_202 & _T_108; // @[AesSbox.scala 41:63]
  wire  _T_236 = _T_200 & _T_88; // @[AesSbox.scala 41:63]
  wire  _T_238 = _T_208 & _T_82; // @[AesSbox.scala 41:63]
  wire  _T_240 = _T_198 & _T_86; // @[AesSbox.scala 41:63]
  wire  _T_242 = _T_196 & _T_112; // @[AesSbox.scala 41:63]
  wire  _T_244 = _T_206 & _T_72; // @[AesSbox.scala 41:63]
  wire  _T_246 = _T_212 & _T_118; // @[AesSbox.scala 41:63]
  wire  _T_248 = _T_204 & _T_100; // @[AesSbox.scala 41:63]
  wire  _T_250 = _T_244 ^ _T_246; // @[AesSbox.scala 40:63]
  wire  _T_252 = _T_222 ^ _T_234; // @[AesSbox.scala 40:63]
  wire  _T_254 = _T_228 ^ _T_250; // @[AesSbox.scala 40:63]
  wire  _T_256 = _T_232 ^ _T_252; // @[AesSbox.scala 40:63]
  wire  _T_258 = _T_218 ^ _T_238; // @[AesSbox.scala 40:63]
  wire  _T_260 = _T_214 ^ _T_220; // @[AesSbox.scala 40:63]
  wire  _T_262 = _T_250 ^ _T_260; // @[AesSbox.scala 40:63]
  wire  _T_264 = _T_216 ^ _T_256; // @[AesSbox.scala 40:63]
  wire  _T_266 = _T_214 ^ _T_226; // @[AesSbox.scala 40:63]
  wire  _T_268 = _T_224 ^ _T_240; // @[AesSbox.scala 40:63]
  wire  _T_270 = _T_230 ^ _T_242; // @[AesSbox.scala 40:63]
  wire  _T_272 = _T_218 ^ _T_264; // @[AesSbox.scala 40:63]
  wire  _T_274 = _T_258 ^ _T_270; // @[AesSbox.scala 40:63]
  wire  _T_276 = _T_236 ^ _T_252; // @[AesSbox.scala 40:63]
  wire  _T_278 = _T_220 ^ _T_226; // @[AesSbox.scala 40:63]
  wire  _T_280 = _T_256 ^ _T_278; // @[AesSbox.scala 40:63]
  wire  _T_282 = _T_248 ^ _T_274; // @[AesSbox.scala 40:63]
  wire  _T_284 = _T_244 ^ _T_266; // @[AesSbox.scala 40:63]
  wire  _T_286 = _T_258 ^ _T_268; // @[AesSbox.scala 40:63]
  wire  _T_287 = _T_254 ^ _T_280; // @[AesSbox.scala 40:63]
  wire  _T_288 = _T_282 ^ _T_284; // @[AesSbox.scala 42:65]
  wire  _T_289 = ~_T_288; // @[AesSbox.scala 42:51]
  wire  _T_291 = _T_224 ^ _T_250; // @[AesSbox.scala 40:63]
  wire  _T_292 = _T_262 ^ _T_264; // @[AesSbox.scala 40:63]
  wire  _T_293 = _T_272 ^ _T_291; // @[AesSbox.scala 40:63]
  wire  _T_295 = _T_222 ^ _T_238; // @[AesSbox.scala 40:63]
  wire  _T_297 = _T_260 ^ _T_276; // @[AesSbox.scala 40:63]
  wire  _T_298 = _T_262 ^ _T_286; // @[AesSbox.scala 42:65]
  wire  _T_299 = ~_T_298; // @[AesSbox.scala 42:51]
  wire  _T_301 = _T_230 ^ _T_268; // @[AesSbox.scala 40:63]
  wire  _T_303 = _T_295 ^ _T_301; // @[AesSbox.scala 40:63]
  wire  _T_305 = _T_222 ^ _T_266; // @[AesSbox.scala 40:63]
  wire  _T_306 = _T_254 ^ _T_303; // @[AesSbox.scala 42:65]
  wire  _T_307 = ~_T_306; // @[AesSbox.scala 42:51]
  wire  _T_309 = _T_274 ^ _T_297; // @[AesSbox.scala 40:63]
  wire  _T_310 = _T_254 ^ _T_309; // @[AesSbox.scala 40:63]
  wire  _T_312 = _T_264 ^ _T_305; // @[AesSbox.scala 40:63]
  wire  _T_313 = _T_254 ^ _T_312; // @[AesSbox.scala 42:65]
  wire  _T_314 = ~_T_313; // @[AesSbox.scala 42:51]
  wire [7:0] _T_321 = {_T_287,_T_314,_T_289,_T_292,_T_293,_T_310,_T_307,_T_299}; // @[Cat.scala 29:58]
  wire  _T_339 = shreg_io_output_0[17] ^ shreg_io_output_0[19]; // @[AesSbox.scala 40:63]
  wire  _T_341 = shreg_io_output_0[20] ^ shreg_io_output_0[23]; // @[AesSbox.scala 40:63]
  wire  _T_343 = shreg_io_output_0[22] ^ shreg_io_output_0[21]; // @[AesSbox.scala 40:63]
  wire  _T_345 = shreg_io_output_0[16] ^ _T_343; // @[AesSbox.scala 40:63]
  wire  _T_347 = _T_339 ^ _T_341; // @[AesSbox.scala 40:63]
  wire  _T_349 = shreg_io_output_0[22] ^ shreg_io_output_0[18]; // @[AesSbox.scala 40:63]
  wire  _T_351 = shreg_io_output_0[23] ^ shreg_io_output_0[17]; // @[AesSbox.scala 40:63]
  wire  _T_353 = _T_339 ^ _T_349; // @[AesSbox.scala 40:63]
  wire  _T_355 = shreg_io_output_0[17] ^ _T_345; // @[AesSbox.scala 40:63]
  wire  _T_357 = shreg_io_output_0[20] ^ _T_345; // @[AesSbox.scala 40:63]
  wire  _T_359 = shreg_io_output_0[16] ^ _T_347; // @[AesSbox.scala 40:63]
  wire  _T_361 = _T_347 ^ _T_349; // @[AesSbox.scala 40:63]
  wire  _T_363 = shreg_io_output_0[21] ^ shreg_io_output_0[18]; // @[AesSbox.scala 40:63]
  wire  _T_365 = _T_343 ^ _T_347; // @[AesSbox.scala 40:63]
  wire  _T_367 = shreg_io_output_0[18] ^ _T_351; // @[AesSbox.scala 40:63]
  wire  _T_369 = shreg_io_output_0[23] ^ shreg_io_output_0[18]; // @[AesSbox.scala 40:63]
  wire  _T_371 = shreg_io_output_0[16] ^ _T_353; // @[AesSbox.scala 40:63]
  wire  _T_373 = shreg_io_output_0[17] ^ shreg_io_output_0[18]; // @[AesSbox.scala 40:63]
  wire  _T_375 = _T_341 ^ _T_373; // @[AesSbox.scala 40:63]
  wire  _T_377 = _T_345 ^ _T_367; // @[AesSbox.scala 40:63]
  wire  _T_379 = _T_339 ^ _T_363; // @[AesSbox.scala 40:63]
  wire  _T_381 = shreg_io_output_0[23] ^ _T_345; // @[AesSbox.scala 40:63]
  wire  _T_383 = _T_379 ^ _T_347; // @[AesSbox.scala 40:63]
  wire  _T_385 = _T_379 ^ _T_351; // @[AesSbox.scala 40:63]
  wire  _T_387 = _T_351 ^ _T_375; // @[AesSbox.scala 40:63]
  wire  _T_389 = _T_369 ^ _T_365; // @[AesSbox.scala 40:63]
  wire  _T_391 = _T_381 ^ _T_371; // @[AesSbox.scala 40:63]
  wire  _T_393 = _T_375 & _T_347; // @[AesSbox.scala 41:63]
  wire  _T_395 = _T_377 & _T_359; // @[AesSbox.scala 41:63]
  wire  _T_397 = _T_361 ^ _T_393; // @[AesSbox.scala 40:63]
  wire  _T_399 = _T_357 & shreg_io_output_0[16]; // @[AesSbox.scala 41:63]
  wire  _T_401 = _T_399 ^ _T_393; // @[AesSbox.scala 40:63]
  wire  _T_403 = _T_351 & _T_379; // @[AesSbox.scala 41:63]
  wire  _T_405 = _T_355 & _T_345; // @[AesSbox.scala 41:63]
  wire  _T_407 = _T_385 ^ _T_403; // @[AesSbox.scala 40:63]
  wire  _T_409 = _T_381 & _T_371; // @[AesSbox.scala 41:63]
  wire  _T_411 = _T_409 ^ _T_403; // @[AesSbox.scala 40:63]
  wire  _T_413 = _T_341 & _T_353; // @[AesSbox.scala 41:63]
  wire  _T_415 = _T_387 & _T_383; // @[AesSbox.scala 41:63]
  wire  _T_417 = _T_415 ^ _T_413; // @[AesSbox.scala 40:63]
  wire  _T_419 = _T_369 & _T_365; // @[AesSbox.scala 41:63]
  wire  _T_421 = _T_419 ^ _T_413; // @[AesSbox.scala 40:63]
  wire  _T_423 = _T_397 ^ _T_395; // @[AesSbox.scala 40:63]
  wire  _T_425 = _T_401 ^ _T_389; // @[AesSbox.scala 40:63]
  wire  _T_427 = _T_407 ^ _T_405; // @[AesSbox.scala 40:63]
  wire  _T_429 = _T_411 ^ _T_421; // @[AesSbox.scala 40:63]
  wire  _T_431 = _T_423 ^ _T_417; // @[AesSbox.scala 40:63]
  wire  _T_433 = _T_425 ^ _T_421; // @[AesSbox.scala 40:63]
  wire  _T_435 = _T_427 ^ _T_417; // @[AesSbox.scala 40:63]
  wire  _T_437 = _T_429 ^ _T_391; // @[AesSbox.scala 40:63]
  wire  _T_439 = _T_435 ^ _T_437; // @[AesSbox.scala 40:63]
  wire  _T_441 = _T_435 & _T_431; // @[AesSbox.scala 41:63]
  wire  _T_443 = _T_433 ^ _T_441; // @[AesSbox.scala 40:63]
  wire  _T_445 = _T_431 ^ _T_433; // @[AesSbox.scala 40:63]
  wire  _T_447 = _T_437 ^ _T_441; // @[AesSbox.scala 40:63]
  wire  _T_449 = _T_447 & _T_445; // @[AesSbox.scala 41:63]
  wire  _T_451 = _T_443 & _T_439; // @[AesSbox.scala 41:63]
  wire  _T_453 = _T_431 & _T_437; // @[AesSbox.scala 41:63]
  wire  _T_455 = _T_445 & _T_453; // @[AesSbox.scala 41:63]
  wire  _T_457 = _T_445 ^ _T_441; // @[AesSbox.scala 40:63]
  wire  _T_459 = _T_433 & _T_435; // @[AesSbox.scala 41:63]
  wire  _T_461 = _T_439 & _T_459; // @[AesSbox.scala 41:63]
  wire  _T_463 = _T_439 ^ _T_441; // @[AesSbox.scala 40:63]
  wire  _T_465 = _T_433 ^ _T_449; // @[AesSbox.scala 40:63]
  wire  _T_467 = _T_455 ^ _T_457; // @[AesSbox.scala 40:63]
  wire  _T_469 = _T_437 ^ _T_451; // @[AesSbox.scala 40:63]
  wire  _T_471 = _T_461 ^ _T_463; // @[AesSbox.scala 40:63]
  wire  _T_473 = _T_467 ^ _T_471; // @[AesSbox.scala 40:63]
  wire  _T_475 = _T_465 ^ _T_469; // @[AesSbox.scala 40:63]
  wire  _T_477 = _T_465 ^ _T_467; // @[AesSbox.scala 40:63]
  wire  _T_479 = _T_469 ^ _T_471; // @[AesSbox.scala 40:63]
  wire  _T_481 = _T_475 ^ _T_473; // @[AesSbox.scala 40:63]
  wire  _T_483 = _T_479 & _T_347; // @[AesSbox.scala 41:63]
  wire  _T_485 = _T_471 & _T_359; // @[AesSbox.scala 41:63]
  wire  _T_487 = _T_469 & shreg_io_output_0[16]; // @[AesSbox.scala 41:63]
  wire  _T_489 = _T_477 & _T_379; // @[AesSbox.scala 41:63]
  wire  _T_491 = _T_467 & _T_345; // @[AesSbox.scala 41:63]
  wire  _T_493 = _T_465 & _T_371; // @[AesSbox.scala 41:63]
  wire  _T_495 = _T_475 & _T_353; // @[AesSbox.scala 41:63]
  wire  _T_497 = _T_481 & _T_383; // @[AesSbox.scala 41:63]
  wire  _T_499 = _T_473 & _T_365; // @[AesSbox.scala 41:63]
  wire  _T_501 = _T_479 & _T_375; // @[AesSbox.scala 41:63]
  wire  _T_503 = _T_471 & _T_377; // @[AesSbox.scala 41:63]
  wire  _T_505 = _T_469 & _T_357; // @[AesSbox.scala 41:63]
  wire  _T_507 = _T_477 & _T_351; // @[AesSbox.scala 41:63]
  wire  _T_509 = _T_467 & _T_355; // @[AesSbox.scala 41:63]
  wire  _T_511 = _T_465 & _T_381; // @[AesSbox.scala 41:63]
  wire  _T_513 = _T_475 & _T_341; // @[AesSbox.scala 41:63]
  wire  _T_515 = _T_481 & _T_387; // @[AesSbox.scala 41:63]
  wire  _T_517 = _T_473 & _T_369; // @[AesSbox.scala 41:63]
  wire  _T_519 = _T_513 ^ _T_515; // @[AesSbox.scala 40:63]
  wire  _T_521 = _T_491 ^ _T_503; // @[AesSbox.scala 40:63]
  wire  _T_523 = _T_497 ^ _T_519; // @[AesSbox.scala 40:63]
  wire  _T_525 = _T_501 ^ _T_521; // @[AesSbox.scala 40:63]
  wire  _T_527 = _T_487 ^ _T_507; // @[AesSbox.scala 40:63]
  wire  _T_529 = _T_483 ^ _T_489; // @[AesSbox.scala 40:63]
  wire  _T_531 = _T_519 ^ _T_529; // @[AesSbox.scala 40:63]
  wire  _T_533 = _T_485 ^ _T_525; // @[AesSbox.scala 40:63]
  wire  _T_535 = _T_483 ^ _T_495; // @[AesSbox.scala 40:63]
  wire  _T_537 = _T_493 ^ _T_509; // @[AesSbox.scala 40:63]
  wire  _T_539 = _T_499 ^ _T_511; // @[AesSbox.scala 40:63]
  wire  _T_541 = _T_487 ^ _T_533; // @[AesSbox.scala 40:63]
  wire  _T_543 = _T_527 ^ _T_539; // @[AesSbox.scala 40:63]
  wire  _T_545 = _T_505 ^ _T_521; // @[AesSbox.scala 40:63]
  wire  _T_547 = _T_489 ^ _T_495; // @[AesSbox.scala 40:63]
  wire  _T_549 = _T_525 ^ _T_547; // @[AesSbox.scala 40:63]
  wire  _T_551 = _T_517 ^ _T_543; // @[AesSbox.scala 40:63]
  wire  _T_553 = _T_513 ^ _T_535; // @[AesSbox.scala 40:63]
  wire  _T_555 = _T_527 ^ _T_537; // @[AesSbox.scala 40:63]
  wire  _T_556 = _T_523 ^ _T_549; // @[AesSbox.scala 40:63]
  wire  _T_557 = _T_551 ^ _T_553; // @[AesSbox.scala 42:65]
  wire  _T_558 = ~_T_557; // @[AesSbox.scala 42:51]
  wire  _T_560 = _T_493 ^ _T_519; // @[AesSbox.scala 40:63]
  wire  _T_561 = _T_531 ^ _T_533; // @[AesSbox.scala 40:63]
  wire  _T_562 = _T_541 ^ _T_560; // @[AesSbox.scala 40:63]
  wire  _T_564 = _T_491 ^ _T_507; // @[AesSbox.scala 40:63]
  wire  _T_566 = _T_529 ^ _T_545; // @[AesSbox.scala 40:63]
  wire  _T_567 = _T_531 ^ _T_555; // @[AesSbox.scala 42:65]
  wire  _T_568 = ~_T_567; // @[AesSbox.scala 42:51]
  wire  _T_570 = _T_499 ^ _T_537; // @[AesSbox.scala 40:63]
  wire  _T_572 = _T_564 ^ _T_570; // @[AesSbox.scala 40:63]
  wire  _T_574 = _T_491 ^ _T_535; // @[AesSbox.scala 40:63]
  wire  _T_575 = _T_523 ^ _T_572; // @[AesSbox.scala 42:65]
  wire  _T_576 = ~_T_575; // @[AesSbox.scala 42:51]
  wire  _T_578 = _T_543 ^ _T_566; // @[AesSbox.scala 40:63]
  wire  _T_579 = _T_523 ^ _T_578; // @[AesSbox.scala 40:63]
  wire  _T_581 = _T_533 ^ _T_574; // @[AesSbox.scala 40:63]
  wire  _T_582 = _T_523 ^ _T_581; // @[AesSbox.scala 42:65]
  wire  _T_583 = ~_T_582; // @[AesSbox.scala 42:51]
  wire [7:0] _T_590 = {_T_556,_T_583,_T_558,_T_561,_T_562,_T_579,_T_576,_T_568}; // @[Cat.scala 29:58]
  wire  _T_608 = shreg_io_output_0[9] ^ shreg_io_output_0[11]; // @[AesSbox.scala 40:63]
  wire  _T_610 = shreg_io_output_0[12] ^ shreg_io_output_0[15]; // @[AesSbox.scala 40:63]
  wire  _T_612 = shreg_io_output_0[14] ^ shreg_io_output_0[13]; // @[AesSbox.scala 40:63]
  wire  _T_614 = shreg_io_output_0[8] ^ _T_612; // @[AesSbox.scala 40:63]
  wire  _T_616 = _T_608 ^ _T_610; // @[AesSbox.scala 40:63]
  wire  _T_618 = shreg_io_output_0[14] ^ shreg_io_output_0[10]; // @[AesSbox.scala 40:63]
  wire  _T_620 = shreg_io_output_0[15] ^ shreg_io_output_0[9]; // @[AesSbox.scala 40:63]
  wire  _T_622 = _T_608 ^ _T_618; // @[AesSbox.scala 40:63]
  wire  _T_624 = shreg_io_output_0[9] ^ _T_614; // @[AesSbox.scala 40:63]
  wire  _T_626 = shreg_io_output_0[12] ^ _T_614; // @[AesSbox.scala 40:63]
  wire  _T_628 = shreg_io_output_0[8] ^ _T_616; // @[AesSbox.scala 40:63]
  wire  _T_630 = _T_616 ^ _T_618; // @[AesSbox.scala 40:63]
  wire  _T_632 = shreg_io_output_0[13] ^ shreg_io_output_0[10]; // @[AesSbox.scala 40:63]
  wire  _T_634 = _T_612 ^ _T_616; // @[AesSbox.scala 40:63]
  wire  _T_636 = shreg_io_output_0[10] ^ _T_620; // @[AesSbox.scala 40:63]
  wire  _T_638 = shreg_io_output_0[15] ^ shreg_io_output_0[10]; // @[AesSbox.scala 40:63]
  wire  _T_640 = shreg_io_output_0[8] ^ _T_622; // @[AesSbox.scala 40:63]
  wire  _T_642 = shreg_io_output_0[9] ^ shreg_io_output_0[10]; // @[AesSbox.scala 40:63]
  wire  _T_644 = _T_610 ^ _T_642; // @[AesSbox.scala 40:63]
  wire  _T_646 = _T_614 ^ _T_636; // @[AesSbox.scala 40:63]
  wire  _T_648 = _T_608 ^ _T_632; // @[AesSbox.scala 40:63]
  wire  _T_650 = shreg_io_output_0[15] ^ _T_614; // @[AesSbox.scala 40:63]
  wire  _T_652 = _T_648 ^ _T_616; // @[AesSbox.scala 40:63]
  wire  _T_654 = _T_648 ^ _T_620; // @[AesSbox.scala 40:63]
  wire  _T_656 = _T_620 ^ _T_644; // @[AesSbox.scala 40:63]
  wire  _T_658 = _T_638 ^ _T_634; // @[AesSbox.scala 40:63]
  wire  _T_660 = _T_650 ^ _T_640; // @[AesSbox.scala 40:63]
  wire  _T_662 = _T_644 & _T_616; // @[AesSbox.scala 41:63]
  wire  _T_664 = _T_646 & _T_628; // @[AesSbox.scala 41:63]
  wire  _T_666 = _T_630 ^ _T_662; // @[AesSbox.scala 40:63]
  wire  _T_668 = _T_626 & shreg_io_output_0[8]; // @[AesSbox.scala 41:63]
  wire  _T_670 = _T_668 ^ _T_662; // @[AesSbox.scala 40:63]
  wire  _T_672 = _T_620 & _T_648; // @[AesSbox.scala 41:63]
  wire  _T_674 = _T_624 & _T_614; // @[AesSbox.scala 41:63]
  wire  _T_676 = _T_654 ^ _T_672; // @[AesSbox.scala 40:63]
  wire  _T_678 = _T_650 & _T_640; // @[AesSbox.scala 41:63]
  wire  _T_680 = _T_678 ^ _T_672; // @[AesSbox.scala 40:63]
  wire  _T_682 = _T_610 & _T_622; // @[AesSbox.scala 41:63]
  wire  _T_684 = _T_656 & _T_652; // @[AesSbox.scala 41:63]
  wire  _T_686 = _T_684 ^ _T_682; // @[AesSbox.scala 40:63]
  wire  _T_688 = _T_638 & _T_634; // @[AesSbox.scala 41:63]
  wire  _T_690 = _T_688 ^ _T_682; // @[AesSbox.scala 40:63]
  wire  _T_692 = _T_666 ^ _T_664; // @[AesSbox.scala 40:63]
  wire  _T_694 = _T_670 ^ _T_658; // @[AesSbox.scala 40:63]
  wire  _T_696 = _T_676 ^ _T_674; // @[AesSbox.scala 40:63]
  wire  _T_698 = _T_680 ^ _T_690; // @[AesSbox.scala 40:63]
  wire  _T_700 = _T_692 ^ _T_686; // @[AesSbox.scala 40:63]
  wire  _T_702 = _T_694 ^ _T_690; // @[AesSbox.scala 40:63]
  wire  _T_704 = _T_696 ^ _T_686; // @[AesSbox.scala 40:63]
  wire  _T_706 = _T_698 ^ _T_660; // @[AesSbox.scala 40:63]
  wire  _T_708 = _T_704 ^ _T_706; // @[AesSbox.scala 40:63]
  wire  _T_710 = _T_704 & _T_700; // @[AesSbox.scala 41:63]
  wire  _T_712 = _T_702 ^ _T_710; // @[AesSbox.scala 40:63]
  wire  _T_714 = _T_700 ^ _T_702; // @[AesSbox.scala 40:63]
  wire  _T_716 = _T_706 ^ _T_710; // @[AesSbox.scala 40:63]
  wire  _T_718 = _T_716 & _T_714; // @[AesSbox.scala 41:63]
  wire  _T_720 = _T_712 & _T_708; // @[AesSbox.scala 41:63]
  wire  _T_722 = _T_700 & _T_706; // @[AesSbox.scala 41:63]
  wire  _T_724 = _T_714 & _T_722; // @[AesSbox.scala 41:63]
  wire  _T_726 = _T_714 ^ _T_710; // @[AesSbox.scala 40:63]
  wire  _T_728 = _T_702 & _T_704; // @[AesSbox.scala 41:63]
  wire  _T_730 = _T_708 & _T_728; // @[AesSbox.scala 41:63]
  wire  _T_732 = _T_708 ^ _T_710; // @[AesSbox.scala 40:63]
  wire  _T_734 = _T_702 ^ _T_718; // @[AesSbox.scala 40:63]
  wire  _T_736 = _T_724 ^ _T_726; // @[AesSbox.scala 40:63]
  wire  _T_738 = _T_706 ^ _T_720; // @[AesSbox.scala 40:63]
  wire  _T_740 = _T_730 ^ _T_732; // @[AesSbox.scala 40:63]
  wire  _T_742 = _T_736 ^ _T_740; // @[AesSbox.scala 40:63]
  wire  _T_744 = _T_734 ^ _T_738; // @[AesSbox.scala 40:63]
  wire  _T_746 = _T_734 ^ _T_736; // @[AesSbox.scala 40:63]
  wire  _T_748 = _T_738 ^ _T_740; // @[AesSbox.scala 40:63]
  wire  _T_750 = _T_744 ^ _T_742; // @[AesSbox.scala 40:63]
  wire  _T_752 = _T_748 & _T_616; // @[AesSbox.scala 41:63]
  wire  _T_754 = _T_740 & _T_628; // @[AesSbox.scala 41:63]
  wire  _T_756 = _T_738 & shreg_io_output_0[8]; // @[AesSbox.scala 41:63]
  wire  _T_758 = _T_746 & _T_648; // @[AesSbox.scala 41:63]
  wire  _T_760 = _T_736 & _T_614; // @[AesSbox.scala 41:63]
  wire  _T_762 = _T_734 & _T_640; // @[AesSbox.scala 41:63]
  wire  _T_764 = _T_744 & _T_622; // @[AesSbox.scala 41:63]
  wire  _T_766 = _T_750 & _T_652; // @[AesSbox.scala 41:63]
  wire  _T_768 = _T_742 & _T_634; // @[AesSbox.scala 41:63]
  wire  _T_770 = _T_748 & _T_644; // @[AesSbox.scala 41:63]
  wire  _T_772 = _T_740 & _T_646; // @[AesSbox.scala 41:63]
  wire  _T_774 = _T_738 & _T_626; // @[AesSbox.scala 41:63]
  wire  _T_776 = _T_746 & _T_620; // @[AesSbox.scala 41:63]
  wire  _T_778 = _T_736 & _T_624; // @[AesSbox.scala 41:63]
  wire  _T_780 = _T_734 & _T_650; // @[AesSbox.scala 41:63]
  wire  _T_782 = _T_744 & _T_610; // @[AesSbox.scala 41:63]
  wire  _T_784 = _T_750 & _T_656; // @[AesSbox.scala 41:63]
  wire  _T_786 = _T_742 & _T_638; // @[AesSbox.scala 41:63]
  wire  _T_788 = _T_782 ^ _T_784; // @[AesSbox.scala 40:63]
  wire  _T_790 = _T_760 ^ _T_772; // @[AesSbox.scala 40:63]
  wire  _T_792 = _T_766 ^ _T_788; // @[AesSbox.scala 40:63]
  wire  _T_794 = _T_770 ^ _T_790; // @[AesSbox.scala 40:63]
  wire  _T_796 = _T_756 ^ _T_776; // @[AesSbox.scala 40:63]
  wire  _T_798 = _T_752 ^ _T_758; // @[AesSbox.scala 40:63]
  wire  _T_800 = _T_788 ^ _T_798; // @[AesSbox.scala 40:63]
  wire  _T_802 = _T_754 ^ _T_794; // @[AesSbox.scala 40:63]
  wire  _T_804 = _T_752 ^ _T_764; // @[AesSbox.scala 40:63]
  wire  _T_806 = _T_762 ^ _T_778; // @[AesSbox.scala 40:63]
  wire  _T_808 = _T_768 ^ _T_780; // @[AesSbox.scala 40:63]
  wire  _T_810 = _T_756 ^ _T_802; // @[AesSbox.scala 40:63]
  wire  _T_812 = _T_796 ^ _T_808; // @[AesSbox.scala 40:63]
  wire  _T_814 = _T_774 ^ _T_790; // @[AesSbox.scala 40:63]
  wire  _T_816 = _T_758 ^ _T_764; // @[AesSbox.scala 40:63]
  wire  _T_818 = _T_794 ^ _T_816; // @[AesSbox.scala 40:63]
  wire  _T_820 = _T_786 ^ _T_812; // @[AesSbox.scala 40:63]
  wire  _T_822 = _T_782 ^ _T_804; // @[AesSbox.scala 40:63]
  wire  _T_824 = _T_796 ^ _T_806; // @[AesSbox.scala 40:63]
  wire  _T_825 = _T_792 ^ _T_818; // @[AesSbox.scala 40:63]
  wire  _T_826 = _T_820 ^ _T_822; // @[AesSbox.scala 42:65]
  wire  _T_827 = ~_T_826; // @[AesSbox.scala 42:51]
  wire  _T_829 = _T_762 ^ _T_788; // @[AesSbox.scala 40:63]
  wire  _T_830 = _T_800 ^ _T_802; // @[AesSbox.scala 40:63]
  wire  _T_831 = _T_810 ^ _T_829; // @[AesSbox.scala 40:63]
  wire  _T_833 = _T_760 ^ _T_776; // @[AesSbox.scala 40:63]
  wire  _T_835 = _T_798 ^ _T_814; // @[AesSbox.scala 40:63]
  wire  _T_836 = _T_800 ^ _T_824; // @[AesSbox.scala 42:65]
  wire  _T_837 = ~_T_836; // @[AesSbox.scala 42:51]
  wire  _T_839 = _T_768 ^ _T_806; // @[AesSbox.scala 40:63]
  wire  _T_841 = _T_833 ^ _T_839; // @[AesSbox.scala 40:63]
  wire  _T_843 = _T_760 ^ _T_804; // @[AesSbox.scala 40:63]
  wire  _T_844 = _T_792 ^ _T_841; // @[AesSbox.scala 42:65]
  wire  _T_845 = ~_T_844; // @[AesSbox.scala 42:51]
  wire  _T_847 = _T_812 ^ _T_835; // @[AesSbox.scala 40:63]
  wire  _T_848 = _T_792 ^ _T_847; // @[AesSbox.scala 40:63]
  wire  _T_850 = _T_802 ^ _T_843; // @[AesSbox.scala 40:63]
  wire  _T_851 = _T_792 ^ _T_850; // @[AesSbox.scala 42:65]
  wire  _T_852 = ~_T_851; // @[AesSbox.scala 42:51]
  wire [7:0] _T_859 = {_T_825,_T_852,_T_827,_T_830,_T_831,_T_848,_T_845,_T_837}; // @[Cat.scala 29:58]
  wire  _T_877 = shreg_io_output_0[1] ^ shreg_io_output_0[3]; // @[AesSbox.scala 40:63]
  wire  _T_879 = shreg_io_output_0[4] ^ shreg_io_output_0[7]; // @[AesSbox.scala 40:63]
  wire  _T_881 = shreg_io_output_0[6] ^ shreg_io_output_0[5]; // @[AesSbox.scala 40:63]
  wire  _T_883 = shreg_io_output_0[0] ^ _T_881; // @[AesSbox.scala 40:63]
  wire  _T_885 = _T_877 ^ _T_879; // @[AesSbox.scala 40:63]
  wire  _T_887 = shreg_io_output_0[6] ^ shreg_io_output_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_889 = shreg_io_output_0[7] ^ shreg_io_output_0[1]; // @[AesSbox.scala 40:63]
  wire  _T_891 = _T_877 ^ _T_887; // @[AesSbox.scala 40:63]
  wire  _T_893 = shreg_io_output_0[1] ^ _T_883; // @[AesSbox.scala 40:63]
  wire  _T_895 = shreg_io_output_0[4] ^ _T_883; // @[AesSbox.scala 40:63]
  wire  _T_897 = shreg_io_output_0[0] ^ _T_885; // @[AesSbox.scala 40:63]
  wire  _T_899 = _T_885 ^ _T_887; // @[AesSbox.scala 40:63]
  wire  _T_901 = shreg_io_output_0[5] ^ shreg_io_output_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_903 = _T_881 ^ _T_885; // @[AesSbox.scala 40:63]
  wire  _T_905 = shreg_io_output_0[2] ^ _T_889; // @[AesSbox.scala 40:63]
  wire  _T_907 = shreg_io_output_0[7] ^ shreg_io_output_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_909 = shreg_io_output_0[0] ^ _T_891; // @[AesSbox.scala 40:63]
  wire  _T_911 = shreg_io_output_0[1] ^ shreg_io_output_0[2]; // @[AesSbox.scala 40:63]
  wire  _T_913 = _T_879 ^ _T_911; // @[AesSbox.scala 40:63]
  wire  _T_915 = _T_883 ^ _T_905; // @[AesSbox.scala 40:63]
  wire  _T_917 = _T_877 ^ _T_901; // @[AesSbox.scala 40:63]
  wire  _T_919 = shreg_io_output_0[7] ^ _T_883; // @[AesSbox.scala 40:63]
  wire  _T_921 = _T_917 ^ _T_885; // @[AesSbox.scala 40:63]
  wire  _T_923 = _T_917 ^ _T_889; // @[AesSbox.scala 40:63]
  wire  _T_925 = _T_889 ^ _T_913; // @[AesSbox.scala 40:63]
  wire  _T_927 = _T_907 ^ _T_903; // @[AesSbox.scala 40:63]
  wire  _T_929 = _T_919 ^ _T_909; // @[AesSbox.scala 40:63]
  wire  _T_931 = _T_913 & _T_885; // @[AesSbox.scala 41:63]
  wire  _T_933 = _T_915 & _T_897; // @[AesSbox.scala 41:63]
  wire  _T_935 = _T_899 ^ _T_931; // @[AesSbox.scala 40:63]
  wire  _T_937 = _T_895 & shreg_io_output_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_939 = _T_937 ^ _T_931; // @[AesSbox.scala 40:63]
  wire  _T_941 = _T_889 & _T_917; // @[AesSbox.scala 41:63]
  wire  _T_943 = _T_893 & _T_883; // @[AesSbox.scala 41:63]
  wire  _T_945 = _T_923 ^ _T_941; // @[AesSbox.scala 40:63]
  wire  _T_947 = _T_919 & _T_909; // @[AesSbox.scala 41:63]
  wire  _T_949 = _T_947 ^ _T_941; // @[AesSbox.scala 40:63]
  wire  _T_951 = _T_879 & _T_891; // @[AesSbox.scala 41:63]
  wire  _T_953 = _T_925 & _T_921; // @[AesSbox.scala 41:63]
  wire  _T_955 = _T_953 ^ _T_951; // @[AesSbox.scala 40:63]
  wire  _T_957 = _T_907 & _T_903; // @[AesSbox.scala 41:63]
  wire  _T_959 = _T_957 ^ _T_951; // @[AesSbox.scala 40:63]
  wire  _T_961 = _T_935 ^ _T_933; // @[AesSbox.scala 40:63]
  wire  _T_963 = _T_939 ^ _T_927; // @[AesSbox.scala 40:63]
  wire  _T_965 = _T_945 ^ _T_943; // @[AesSbox.scala 40:63]
  wire  _T_967 = _T_949 ^ _T_959; // @[AesSbox.scala 40:63]
  wire  _T_969 = _T_961 ^ _T_955; // @[AesSbox.scala 40:63]
  wire  _T_971 = _T_963 ^ _T_959; // @[AesSbox.scala 40:63]
  wire  _T_973 = _T_965 ^ _T_955; // @[AesSbox.scala 40:63]
  wire  _T_975 = _T_967 ^ _T_929; // @[AesSbox.scala 40:63]
  wire  _T_977 = _T_973 ^ _T_975; // @[AesSbox.scala 40:63]
  wire  _T_979 = _T_973 & _T_969; // @[AesSbox.scala 41:63]
  wire  _T_981 = _T_971 ^ _T_979; // @[AesSbox.scala 40:63]
  wire  _T_983 = _T_969 ^ _T_971; // @[AesSbox.scala 40:63]
  wire  _T_985 = _T_975 ^ _T_979; // @[AesSbox.scala 40:63]
  wire  _T_987 = _T_985 & _T_983; // @[AesSbox.scala 41:63]
  wire  _T_989 = _T_981 & _T_977; // @[AesSbox.scala 41:63]
  wire  _T_991 = _T_969 & _T_975; // @[AesSbox.scala 41:63]
  wire  _T_993 = _T_983 & _T_991; // @[AesSbox.scala 41:63]
  wire  _T_995 = _T_983 ^ _T_979; // @[AesSbox.scala 40:63]
  wire  _T_997 = _T_971 & _T_973; // @[AesSbox.scala 41:63]
  wire  _T_999 = _T_977 & _T_997; // @[AesSbox.scala 41:63]
  wire  _T_1001 = _T_977 ^ _T_979; // @[AesSbox.scala 40:63]
  wire  _T_1003 = _T_971 ^ _T_987; // @[AesSbox.scala 40:63]
  wire  _T_1005 = _T_993 ^ _T_995; // @[AesSbox.scala 40:63]
  wire  _T_1007 = _T_975 ^ _T_989; // @[AesSbox.scala 40:63]
  wire  _T_1009 = _T_999 ^ _T_1001; // @[AesSbox.scala 40:63]
  wire  _T_1011 = _T_1005 ^ _T_1009; // @[AesSbox.scala 40:63]
  wire  _T_1013 = _T_1003 ^ _T_1007; // @[AesSbox.scala 40:63]
  wire  _T_1015 = _T_1003 ^ _T_1005; // @[AesSbox.scala 40:63]
  wire  _T_1017 = _T_1007 ^ _T_1009; // @[AesSbox.scala 40:63]
  wire  _T_1019 = _T_1013 ^ _T_1011; // @[AesSbox.scala 40:63]
  wire  _T_1021 = _T_1017 & _T_885; // @[AesSbox.scala 41:63]
  wire  _T_1023 = _T_1009 & _T_897; // @[AesSbox.scala 41:63]
  wire  _T_1025 = _T_1007 & shreg_io_output_0[0]; // @[AesSbox.scala 41:63]
  wire  _T_1027 = _T_1015 & _T_917; // @[AesSbox.scala 41:63]
  wire  _T_1029 = _T_1005 & _T_883; // @[AesSbox.scala 41:63]
  wire  _T_1031 = _T_1003 & _T_909; // @[AesSbox.scala 41:63]
  wire  _T_1033 = _T_1013 & _T_891; // @[AesSbox.scala 41:63]
  wire  _T_1035 = _T_1019 & _T_921; // @[AesSbox.scala 41:63]
  wire  _T_1037 = _T_1011 & _T_903; // @[AesSbox.scala 41:63]
  wire  _T_1039 = _T_1017 & _T_913; // @[AesSbox.scala 41:63]
  wire  _T_1041 = _T_1009 & _T_915; // @[AesSbox.scala 41:63]
  wire  _T_1043 = _T_1007 & _T_895; // @[AesSbox.scala 41:63]
  wire  _T_1045 = _T_1015 & _T_889; // @[AesSbox.scala 41:63]
  wire  _T_1047 = _T_1005 & _T_893; // @[AesSbox.scala 41:63]
  wire  _T_1049 = _T_1003 & _T_919; // @[AesSbox.scala 41:63]
  wire  _T_1051 = _T_1013 & _T_879; // @[AesSbox.scala 41:63]
  wire  _T_1053 = _T_1019 & _T_925; // @[AesSbox.scala 41:63]
  wire  _T_1055 = _T_1011 & _T_907; // @[AesSbox.scala 41:63]
  wire  _T_1057 = _T_1051 ^ _T_1053; // @[AesSbox.scala 40:63]
  wire  _T_1059 = _T_1029 ^ _T_1041; // @[AesSbox.scala 40:63]
  wire  _T_1061 = _T_1035 ^ _T_1057; // @[AesSbox.scala 40:63]
  wire  _T_1063 = _T_1039 ^ _T_1059; // @[AesSbox.scala 40:63]
  wire  _T_1065 = _T_1025 ^ _T_1045; // @[AesSbox.scala 40:63]
  wire  _T_1067 = _T_1021 ^ _T_1027; // @[AesSbox.scala 40:63]
  wire  _T_1069 = _T_1057 ^ _T_1067; // @[AesSbox.scala 40:63]
  wire  _T_1071 = _T_1023 ^ _T_1063; // @[AesSbox.scala 40:63]
  wire  _T_1073 = _T_1021 ^ _T_1033; // @[AesSbox.scala 40:63]
  wire  _T_1075 = _T_1031 ^ _T_1047; // @[AesSbox.scala 40:63]
  wire  _T_1077 = _T_1037 ^ _T_1049; // @[AesSbox.scala 40:63]
  wire  _T_1079 = _T_1025 ^ _T_1071; // @[AesSbox.scala 40:63]
  wire  _T_1081 = _T_1065 ^ _T_1077; // @[AesSbox.scala 40:63]
  wire  _T_1083 = _T_1043 ^ _T_1059; // @[AesSbox.scala 40:63]
  wire  _T_1085 = _T_1027 ^ _T_1033; // @[AesSbox.scala 40:63]
  wire  _T_1087 = _T_1063 ^ _T_1085; // @[AesSbox.scala 40:63]
  wire  _T_1089 = _T_1055 ^ _T_1081; // @[AesSbox.scala 40:63]
  wire  _T_1091 = _T_1051 ^ _T_1073; // @[AesSbox.scala 40:63]
  wire  _T_1093 = _T_1065 ^ _T_1075; // @[AesSbox.scala 40:63]
  wire  _T_1094 = _T_1061 ^ _T_1087; // @[AesSbox.scala 40:63]
  wire  _T_1095 = _T_1089 ^ _T_1091; // @[AesSbox.scala 42:65]
  wire  _T_1096 = ~_T_1095; // @[AesSbox.scala 42:51]
  wire  _T_1098 = _T_1031 ^ _T_1057; // @[AesSbox.scala 40:63]
  wire  _T_1099 = _T_1069 ^ _T_1071; // @[AesSbox.scala 40:63]
  wire  _T_1100 = _T_1079 ^ _T_1098; // @[AesSbox.scala 40:63]
  wire  _T_1102 = _T_1029 ^ _T_1045; // @[AesSbox.scala 40:63]
  wire  _T_1104 = _T_1067 ^ _T_1083; // @[AesSbox.scala 40:63]
  wire  _T_1105 = _T_1069 ^ _T_1093; // @[AesSbox.scala 42:65]
  wire  _T_1106 = ~_T_1105; // @[AesSbox.scala 42:51]
  wire  _T_1108 = _T_1037 ^ _T_1075; // @[AesSbox.scala 40:63]
  wire  _T_1110 = _T_1102 ^ _T_1108; // @[AesSbox.scala 40:63]
  wire  _T_1112 = _T_1029 ^ _T_1073; // @[AesSbox.scala 40:63]
  wire  _T_1113 = _T_1061 ^ _T_1110; // @[AesSbox.scala 42:65]
  wire  _T_1114 = ~_T_1113; // @[AesSbox.scala 42:51]
  wire  _T_1116 = _T_1081 ^ _T_1104; // @[AesSbox.scala 40:63]
  wire  _T_1117 = _T_1061 ^ _T_1116; // @[AesSbox.scala 40:63]
  wire  _T_1119 = _T_1071 ^ _T_1112; // @[AesSbox.scala 40:63]
  wire  _T_1120 = _T_1061 ^ _T_1119; // @[AesSbox.scala 42:65]
  wire  _T_1121 = ~_T_1120; // @[AesSbox.scala 42:51]
  wire [7:0] _T_1128 = {_T_1094,_T_1121,_T_1096,_T_1099,_T_1100,_T_1117,_T_1114,_T_1106}; // @[Cat.scala 29:58]
  wire [7:0] _T_1129_0_0 = io_aes256 ? shreg_io_output_1[127:120] : shreg_io_output_0[127:120]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_0_1 = io_aes256 ? shreg_io_output_1[119:112] : shreg_io_output_0[119:112]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_0_2 = io_aes256 ? shreg_io_output_1[111:104] : shreg_io_output_0[111:104]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_0_3 = io_aes256 ? shreg_io_output_1[103:96] : shreg_io_output_0[103:96]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_1_0 = io_aes256 ? shreg_io_output_1[95:88] : shreg_io_output_0[95:88]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_1_1 = io_aes256 ? shreg_io_output_1[87:80] : shreg_io_output_0[87:80]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_1_2 = io_aes256 ? shreg_io_output_1[79:72] : shreg_io_output_0[79:72]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_1_3 = io_aes256 ? shreg_io_output_1[71:64] : shreg_io_output_0[71:64]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_2_0 = io_aes256 ? shreg_io_output_1[63:56] : shreg_io_output_0[63:56]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_2_1 = io_aes256 ? shreg_io_output_1[55:48] : shreg_io_output_0[55:48]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_2_2 = io_aes256 ? shreg_io_output_1[47:40] : shreg_io_output_0[47:40]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_2_3 = io_aes256 ? shreg_io_output_1[39:32] : shreg_io_output_0[39:32]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_3_0 = io_aes256 ? shreg_io_output_1[31:24] : shreg_io_output_0[31:24]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_3_1 = io_aes256 ? shreg_io_output_1[23:16] : shreg_io_output_0[23:16]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_3_2 = io_aes256 ? shreg_io_output_1[15:8] : shreg_io_output_0[15:8]; // @[AesComponents.scala 121:29]
  wire [7:0] _T_1129_3_3 = io_aes256 ? shreg_io_output_1[7:0] : shreg_io_output_0[7:0]; // @[AesComponents.scala 121:29]
  wire [4:0] _T_1133 = keyInd[5:1] + 5'h1; // @[AesComponents.scala 123:78]
  wire [7:0] _GEN_6 = 4'h1 == _T_1133[3:0] ? 8'h1 : 8'h0; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_7 = 4'h2 == _T_1133[3:0] ? 8'h2 : _GEN_6; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_8 = 4'h3 == _T_1133[3:0] ? 8'h4 : _GEN_7; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_9 = 4'h4 == _T_1133[3:0] ? 8'h8 : _GEN_8; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_10 = 4'h5 == _T_1133[3:0] ? 8'h10 : _GEN_9; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_11 = 4'h6 == _T_1133[3:0] ? 8'h20 : _GEN_10; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_12 = 4'h7 == _T_1133[3:0] ? 8'h40 : _GEN_11; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_13 = 4'h8 == _T_1133[3:0] ? 8'h80 : _GEN_12; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_14 = 4'h9 == _T_1133[3:0] ? 8'h1b : _GEN_13; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_15 = 4'ha == _T_1133[3:0] ? 8'h36 : _GEN_14; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_16 = 4'hb == _T_1133[3:0] ? 8'h6c : _GEN_15; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_17 = 4'hc == _T_1133[3:0] ? 8'hd8 : _GEN_16; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_18 = 4'hd == _T_1133[3:0] ? 8'hab : _GEN_17; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_19 = 4'he == _T_1133[3:0] ? 8'h4d : _GEN_18; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_20 = 4'hf == _T_1133[3:0] ? 8'h9a : _GEN_19; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_22 = 4'h1 == keyInd[3:0] ? 8'h1 : 8'h0; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_23 = 4'h2 == keyInd[3:0] ? 8'h2 : _GEN_22; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_24 = 4'h3 == keyInd[3:0] ? 8'h4 : _GEN_23; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_25 = 4'h4 == keyInd[3:0] ? 8'h8 : _GEN_24; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_26 = 4'h5 == keyInd[3:0] ? 8'h10 : _GEN_25; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_27 = 4'h6 == keyInd[3:0] ? 8'h20 : _GEN_26; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_28 = 4'h7 == keyInd[3:0] ? 8'h40 : _GEN_27; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_29 = 4'h8 == keyInd[3:0] ? 8'h80 : _GEN_28; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_30 = 4'h9 == keyInd[3:0] ? 8'h1b : _GEN_29; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_31 = 4'ha == keyInd[3:0] ? 8'h36 : _GEN_30; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_32 = 4'hb == keyInd[3:0] ? 8'h6c : _GEN_31; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_33 = 4'hc == keyInd[3:0] ? 8'hd8 : _GEN_32; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_34 = 4'hd == keyInd[3:0] ? 8'hab : _GEN_33; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_35 = 4'he == keyInd[3:0] ? 8'h4d : _GEN_34; // @[AesComponents.scala 123:29]
  wire [7:0] _GEN_36 = 4'hf == keyInd[3:0] ? 8'h9a : _GEN_35; // @[AesComponents.scala 123:29]
  wire [7:0] _T_1137 = io_aes256 ? _GEN_20 : _GEN_36; // @[AesComponents.scala 123:29]
  wire [7:0] _T_1138 = _T_52 ? _T_321 : _T_590; // @[AesComponents.scala 125:42]
  wire [7:0] _T_1139 = _T_1129_0_0 ^ _T_1138; // @[AesComponents.scala 125:37]
  wire [7:0] _T_1140 = _T_52 ? 8'h0 : _T_1137; // @[AesComponents.scala 125:67]
  wire [7:0] _T_1141 = _T_1139 ^ _T_1140; // @[AesComponents.scala 125:62]
  wire [7:0] _T_1142 = _T_52 ? _T_590 : _T_859; // @[AesComponents.scala 126:42]
  wire [7:0] _T_1143 = _T_1129_0_1 ^ _T_1142; // @[AesComponents.scala 126:37]
  wire [7:0] _T_1144 = _T_52 ? _T_859 : _T_1128; // @[AesComponents.scala 127:42]
  wire [7:0] _T_1145 = _T_1129_0_2 ^ _T_1144; // @[AesComponents.scala 127:37]
  wire [7:0] _T_1146 = _T_52 ? _T_1128 : _T_321; // @[AesComponents.scala 128:42]
  wire [7:0] _T_1147 = _T_1129_0_3 ^ _T_1146; // @[AesComponents.scala 128:37]
  wire [7:0] _T_1149 = _T_1129_1_0 ^ _T_1141; // @[AesComponents.scala 131:37]
  wire [7:0] _T_1150 = _T_1129_1_1 ^ _T_1143; // @[AesComponents.scala 132:37]
  wire [7:0] _T_1151 = _T_1129_1_2 ^ _T_1145; // @[AesComponents.scala 133:37]
  wire [7:0] _T_1152 = _T_1129_1_3 ^ _T_1147; // @[AesComponents.scala 134:37]
  wire [7:0] _T_1154 = _T_1129_2_0 ^ _T_1149; // @[AesComponents.scala 137:37]
  wire [7:0] _T_1155 = _T_1129_2_1 ^ _T_1150; // @[AesComponents.scala 138:37]
  wire [7:0] _T_1156 = _T_1129_2_2 ^ _T_1151; // @[AesComponents.scala 139:37]
  wire [7:0] _T_1157 = _T_1129_2_3 ^ _T_1152; // @[AesComponents.scala 140:37]
  wire [7:0] _T_1159 = _T_1129_3_0 ^ _T_1154; // @[AesComponents.scala 143:37]
  wire [7:0] _T_1160 = _T_1129_3_1 ^ _T_1155; // @[AesComponents.scala 144:37]
  wire [7:0] _T_1161 = _T_1129_3_2 ^ _T_1156; // @[AesComponents.scala 145:37]
  wire [7:0] _T_1162 = _T_1129_3_3 ^ _T_1157; // @[AesComponents.scala 146:37]
  wire [63:0] _T_1170 = {_T_1154,_T_1155,_T_1156,_T_1157,_T_1159,_T_1160,_T_1161,_T_1162}; // @[Cat.scala 29:58]
  wire [127:0] _T_1178 = {_T_1141,_T_1143,_T_1145,_T_1147,_T_1149,_T_1150,_T_1151,_T_1152,_T_1170}; // @[Cat.scala 29:58]
  wire  _GEN_39 = keyUpdate | _T; // @[AesCombined.scala 71:22]
  wire  _T_1494 = ~keyUpdate; // @[AesCombined.scala 91:36]
  wire  _T_1495 = enc_io_ready & _T_1494; // @[AesCombined.scala 91:33]
  wire  _T_1496 = ~io_keyValid; // @[AesCombined.scala 91:50]
  wire  _T_1499 = dec_io_ready & _T_1494; // @[AesCombined.scala 104:33]
  wire  _T_1504 = enc_io_shift | dec_io_shift; // @[AesCombined.scala 111:24]
  ShiftRegister shreg ( // @[AesCombined.scala 55:23]
    .clock(shreg_clock),
    .io_input(shreg_io_input),
    .io_enable(shreg_io_enable),
    .io_rev(shreg_io_rev),
    .io_cyc(shreg_io_cyc),
    .io_tap(shreg_io_tap),
    .io_output_0(shreg_io_output_0),
    .io_output_1(shreg_io_output_1),
    .io_output_2(shreg_io_output_2),
    .io_output_3(shreg_io_output_3),
    .io_output_4(shreg_io_output_4),
    .io_output_5(shreg_io_output_5),
    .io_output_6(shreg_io_output_6),
    .io_output_7(shreg_io_output_7),
    .io_output_8(shreg_io_output_8),
    .io_output_9(shreg_io_output_9),
    .io_output_10(shreg_io_output_10),
    .io_output_11(shreg_io_output_11),
    .io_output_12(shreg_io_output_12),
    .io_output_13(shreg_io_output_13),
    .io_output_14(shreg_io_output_14)
  );
  AesEncrypt enc ( // @[AesCombined.scala 84:21]
    .clock(enc_clock),
    .reset(enc_reset),
    .io_dataIn(enc_io_dataIn),
    .io_ivIn(enc_io_ivIn),
    .io_dataValid(enc_io_dataValid),
    .io_keys_0_0_0(enc_io_keys_0_0_0),
    .io_keys_0_0_1(enc_io_keys_0_0_1),
    .io_keys_0_0_2(enc_io_keys_0_0_2),
    .io_keys_0_0_3(enc_io_keys_0_0_3),
    .io_keys_0_1_0(enc_io_keys_0_1_0),
    .io_keys_0_1_1(enc_io_keys_0_1_1),
    .io_keys_0_1_2(enc_io_keys_0_1_2),
    .io_keys_0_1_3(enc_io_keys_0_1_3),
    .io_keys_0_2_0(enc_io_keys_0_2_0),
    .io_keys_0_2_1(enc_io_keys_0_2_1),
    .io_keys_0_2_2(enc_io_keys_0_2_2),
    .io_keys_0_2_3(enc_io_keys_0_2_3),
    .io_keys_0_3_0(enc_io_keys_0_3_0),
    .io_keys_0_3_1(enc_io_keys_0_3_1),
    .io_keys_0_3_2(enc_io_keys_0_3_2),
    .io_keys_0_3_3(enc_io_keys_0_3_3),
    .io_aes256(enc_io_aes256),
    .io_shiftCyc(enc_io_shiftCyc),
    .io_shift(enc_io_shift),
    .io_ready(enc_io_ready),
    .io_dataOut(enc_io_dataOut),
    .io_ivOut(enc_io_ivOut),
    .io_outputValid(enc_io_outputValid)
  );
  AesDecrypt dec ( // @[AesCombined.scala 97:21]
    .clock(dec_clock),
    .reset(dec_reset),
    .io_dataIn(dec_io_dataIn),
    .io_ivIn(dec_io_ivIn),
    .io_dataValid(dec_io_dataValid),
    .io_keys_0_0_0(dec_io_keys_0_0_0),
    .io_keys_0_0_1(dec_io_keys_0_0_1),
    .io_keys_0_0_2(dec_io_keys_0_0_2),
    .io_keys_0_0_3(dec_io_keys_0_0_3),
    .io_keys_0_1_0(dec_io_keys_0_1_0),
    .io_keys_0_1_1(dec_io_keys_0_1_1),
    .io_keys_0_1_2(dec_io_keys_0_1_2),
    .io_keys_0_1_3(dec_io_keys_0_1_3),
    .io_keys_0_2_0(dec_io_keys_0_2_0),
    .io_keys_0_2_1(dec_io_keys_0_2_1),
    .io_keys_0_2_2(dec_io_keys_0_2_2),
    .io_keys_0_2_3(dec_io_keys_0_2_3),
    .io_keys_0_3_0(dec_io_keys_0_3_0),
    .io_keys_0_3_1(dec_io_keys_0_3_1),
    .io_keys_0_3_2(dec_io_keys_0_3_2),
    .io_keys_0_3_3(dec_io_keys_0_3_3),
    .io_keys_1_0_0(dec_io_keys_1_0_0),
    .io_keys_1_0_1(dec_io_keys_1_0_1),
    .io_keys_1_0_2(dec_io_keys_1_0_2),
    .io_keys_1_0_3(dec_io_keys_1_0_3),
    .io_keys_1_1_0(dec_io_keys_1_1_0),
    .io_keys_1_1_1(dec_io_keys_1_1_1),
    .io_keys_1_1_2(dec_io_keys_1_1_2),
    .io_keys_1_1_3(dec_io_keys_1_1_3),
    .io_keys_1_2_0(dec_io_keys_1_2_0),
    .io_keys_1_2_1(dec_io_keys_1_2_1),
    .io_keys_1_2_2(dec_io_keys_1_2_2),
    .io_keys_1_2_3(dec_io_keys_1_2_3),
    .io_keys_1_3_0(dec_io_keys_1_3_0),
    .io_keys_1_3_1(dec_io_keys_1_3_1),
    .io_keys_1_3_2(dec_io_keys_1_3_2),
    .io_keys_1_3_3(dec_io_keys_1_3_3),
    .io_keys_2_0_0(dec_io_keys_2_0_0),
    .io_keys_2_0_1(dec_io_keys_2_0_1),
    .io_keys_2_0_2(dec_io_keys_2_0_2),
    .io_keys_2_0_3(dec_io_keys_2_0_3),
    .io_keys_2_1_0(dec_io_keys_2_1_0),
    .io_keys_2_1_1(dec_io_keys_2_1_1),
    .io_keys_2_1_2(dec_io_keys_2_1_2),
    .io_keys_2_1_3(dec_io_keys_2_1_3),
    .io_keys_2_2_0(dec_io_keys_2_2_0),
    .io_keys_2_2_1(dec_io_keys_2_2_1),
    .io_keys_2_2_2(dec_io_keys_2_2_2),
    .io_keys_2_2_3(dec_io_keys_2_2_3),
    .io_keys_2_3_0(dec_io_keys_2_3_0),
    .io_keys_2_3_1(dec_io_keys_2_3_1),
    .io_keys_2_3_2(dec_io_keys_2_3_2),
    .io_keys_2_3_3(dec_io_keys_2_3_3),
    .io_keys_3_0_0(dec_io_keys_3_0_0),
    .io_keys_3_0_1(dec_io_keys_3_0_1),
    .io_keys_3_0_2(dec_io_keys_3_0_2),
    .io_keys_3_0_3(dec_io_keys_3_0_3),
    .io_keys_3_1_0(dec_io_keys_3_1_0),
    .io_keys_3_1_1(dec_io_keys_3_1_1),
    .io_keys_3_1_2(dec_io_keys_3_1_2),
    .io_keys_3_1_3(dec_io_keys_3_1_3),
    .io_keys_3_2_0(dec_io_keys_3_2_0),
    .io_keys_3_2_1(dec_io_keys_3_2_1),
    .io_keys_3_2_2(dec_io_keys_3_2_2),
    .io_keys_3_2_3(dec_io_keys_3_2_3),
    .io_keys_3_3_0(dec_io_keys_3_3_0),
    .io_keys_3_3_1(dec_io_keys_3_3_1),
    .io_keys_3_3_2(dec_io_keys_3_3_2),
    .io_keys_3_3_3(dec_io_keys_3_3_3),
    .io_keys_4_0_0(dec_io_keys_4_0_0),
    .io_keys_4_0_1(dec_io_keys_4_0_1),
    .io_keys_4_0_2(dec_io_keys_4_0_2),
    .io_keys_4_0_3(dec_io_keys_4_0_3),
    .io_keys_4_1_0(dec_io_keys_4_1_0),
    .io_keys_4_1_1(dec_io_keys_4_1_1),
    .io_keys_4_1_2(dec_io_keys_4_1_2),
    .io_keys_4_1_3(dec_io_keys_4_1_3),
    .io_keys_4_2_0(dec_io_keys_4_2_0),
    .io_keys_4_2_1(dec_io_keys_4_2_1),
    .io_keys_4_2_2(dec_io_keys_4_2_2),
    .io_keys_4_2_3(dec_io_keys_4_2_3),
    .io_keys_4_3_0(dec_io_keys_4_3_0),
    .io_keys_4_3_1(dec_io_keys_4_3_1),
    .io_keys_4_3_2(dec_io_keys_4_3_2),
    .io_keys_4_3_3(dec_io_keys_4_3_3),
    .io_keys_5_0_0(dec_io_keys_5_0_0),
    .io_keys_5_0_1(dec_io_keys_5_0_1),
    .io_keys_5_0_2(dec_io_keys_5_0_2),
    .io_keys_5_0_3(dec_io_keys_5_0_3),
    .io_keys_5_1_0(dec_io_keys_5_1_0),
    .io_keys_5_1_1(dec_io_keys_5_1_1),
    .io_keys_5_1_2(dec_io_keys_5_1_2),
    .io_keys_5_1_3(dec_io_keys_5_1_3),
    .io_keys_5_2_0(dec_io_keys_5_2_0),
    .io_keys_5_2_1(dec_io_keys_5_2_1),
    .io_keys_5_2_2(dec_io_keys_5_2_2),
    .io_keys_5_2_3(dec_io_keys_5_2_3),
    .io_keys_5_3_0(dec_io_keys_5_3_0),
    .io_keys_5_3_1(dec_io_keys_5_3_1),
    .io_keys_5_3_2(dec_io_keys_5_3_2),
    .io_keys_5_3_3(dec_io_keys_5_3_3),
    .io_keys_6_0_0(dec_io_keys_6_0_0),
    .io_keys_6_0_1(dec_io_keys_6_0_1),
    .io_keys_6_0_2(dec_io_keys_6_0_2),
    .io_keys_6_0_3(dec_io_keys_6_0_3),
    .io_keys_6_1_0(dec_io_keys_6_1_0),
    .io_keys_6_1_1(dec_io_keys_6_1_1),
    .io_keys_6_1_2(dec_io_keys_6_1_2),
    .io_keys_6_1_3(dec_io_keys_6_1_3),
    .io_keys_6_2_0(dec_io_keys_6_2_0),
    .io_keys_6_2_1(dec_io_keys_6_2_1),
    .io_keys_6_2_2(dec_io_keys_6_2_2),
    .io_keys_6_2_3(dec_io_keys_6_2_3),
    .io_keys_6_3_0(dec_io_keys_6_3_0),
    .io_keys_6_3_1(dec_io_keys_6_3_1),
    .io_keys_6_3_2(dec_io_keys_6_3_2),
    .io_keys_6_3_3(dec_io_keys_6_3_3),
    .io_keys_7_0_0(dec_io_keys_7_0_0),
    .io_keys_7_0_1(dec_io_keys_7_0_1),
    .io_keys_7_0_2(dec_io_keys_7_0_2),
    .io_keys_7_0_3(dec_io_keys_7_0_3),
    .io_keys_7_1_0(dec_io_keys_7_1_0),
    .io_keys_7_1_1(dec_io_keys_7_1_1),
    .io_keys_7_1_2(dec_io_keys_7_1_2),
    .io_keys_7_1_3(dec_io_keys_7_1_3),
    .io_keys_7_2_0(dec_io_keys_7_2_0),
    .io_keys_7_2_1(dec_io_keys_7_2_1),
    .io_keys_7_2_2(dec_io_keys_7_2_2),
    .io_keys_7_2_3(dec_io_keys_7_2_3),
    .io_keys_7_3_0(dec_io_keys_7_3_0),
    .io_keys_7_3_1(dec_io_keys_7_3_1),
    .io_keys_7_3_2(dec_io_keys_7_3_2),
    .io_keys_7_3_3(dec_io_keys_7_3_3),
    .io_keys_8_0_0(dec_io_keys_8_0_0),
    .io_keys_8_0_1(dec_io_keys_8_0_1),
    .io_keys_8_0_2(dec_io_keys_8_0_2),
    .io_keys_8_0_3(dec_io_keys_8_0_3),
    .io_keys_8_1_0(dec_io_keys_8_1_0),
    .io_keys_8_1_1(dec_io_keys_8_1_1),
    .io_keys_8_1_2(dec_io_keys_8_1_2),
    .io_keys_8_1_3(dec_io_keys_8_1_3),
    .io_keys_8_2_0(dec_io_keys_8_2_0),
    .io_keys_8_2_1(dec_io_keys_8_2_1),
    .io_keys_8_2_2(dec_io_keys_8_2_2),
    .io_keys_8_2_3(dec_io_keys_8_2_3),
    .io_keys_8_3_0(dec_io_keys_8_3_0),
    .io_keys_8_3_1(dec_io_keys_8_3_1),
    .io_keys_8_3_2(dec_io_keys_8_3_2),
    .io_keys_8_3_3(dec_io_keys_8_3_3),
    .io_keys_9_0_0(dec_io_keys_9_0_0),
    .io_keys_9_0_1(dec_io_keys_9_0_1),
    .io_keys_9_0_2(dec_io_keys_9_0_2),
    .io_keys_9_0_3(dec_io_keys_9_0_3),
    .io_keys_9_1_0(dec_io_keys_9_1_0),
    .io_keys_9_1_1(dec_io_keys_9_1_1),
    .io_keys_9_1_2(dec_io_keys_9_1_2),
    .io_keys_9_1_3(dec_io_keys_9_1_3),
    .io_keys_9_2_0(dec_io_keys_9_2_0),
    .io_keys_9_2_1(dec_io_keys_9_2_1),
    .io_keys_9_2_2(dec_io_keys_9_2_2),
    .io_keys_9_2_3(dec_io_keys_9_2_3),
    .io_keys_9_3_0(dec_io_keys_9_3_0),
    .io_keys_9_3_1(dec_io_keys_9_3_1),
    .io_keys_9_3_2(dec_io_keys_9_3_2),
    .io_keys_9_3_3(dec_io_keys_9_3_3),
    .io_keys_10_0_0(dec_io_keys_10_0_0),
    .io_keys_10_0_1(dec_io_keys_10_0_1),
    .io_keys_10_0_2(dec_io_keys_10_0_2),
    .io_keys_10_0_3(dec_io_keys_10_0_3),
    .io_keys_10_1_0(dec_io_keys_10_1_0),
    .io_keys_10_1_1(dec_io_keys_10_1_1),
    .io_keys_10_1_2(dec_io_keys_10_1_2),
    .io_keys_10_1_3(dec_io_keys_10_1_3),
    .io_keys_10_2_0(dec_io_keys_10_2_0),
    .io_keys_10_2_1(dec_io_keys_10_2_1),
    .io_keys_10_2_2(dec_io_keys_10_2_2),
    .io_keys_10_2_3(dec_io_keys_10_2_3),
    .io_keys_10_3_0(dec_io_keys_10_3_0),
    .io_keys_10_3_1(dec_io_keys_10_3_1),
    .io_keys_10_3_2(dec_io_keys_10_3_2),
    .io_keys_10_3_3(dec_io_keys_10_3_3),
    .io_keys_11_0_0(dec_io_keys_11_0_0),
    .io_keys_11_0_1(dec_io_keys_11_0_1),
    .io_keys_11_0_2(dec_io_keys_11_0_2),
    .io_keys_11_0_3(dec_io_keys_11_0_3),
    .io_keys_11_1_0(dec_io_keys_11_1_0),
    .io_keys_11_1_1(dec_io_keys_11_1_1),
    .io_keys_11_1_2(dec_io_keys_11_1_2),
    .io_keys_11_1_3(dec_io_keys_11_1_3),
    .io_keys_11_2_0(dec_io_keys_11_2_0),
    .io_keys_11_2_1(dec_io_keys_11_2_1),
    .io_keys_11_2_2(dec_io_keys_11_2_2),
    .io_keys_11_2_3(dec_io_keys_11_2_3),
    .io_keys_11_3_0(dec_io_keys_11_3_0),
    .io_keys_11_3_1(dec_io_keys_11_3_1),
    .io_keys_11_3_2(dec_io_keys_11_3_2),
    .io_keys_11_3_3(dec_io_keys_11_3_3),
    .io_keys_12_0_0(dec_io_keys_12_0_0),
    .io_keys_12_0_1(dec_io_keys_12_0_1),
    .io_keys_12_0_2(dec_io_keys_12_0_2),
    .io_keys_12_0_3(dec_io_keys_12_0_3),
    .io_keys_12_1_0(dec_io_keys_12_1_0),
    .io_keys_12_1_1(dec_io_keys_12_1_1),
    .io_keys_12_1_2(dec_io_keys_12_1_2),
    .io_keys_12_1_3(dec_io_keys_12_1_3),
    .io_keys_12_2_0(dec_io_keys_12_2_0),
    .io_keys_12_2_1(dec_io_keys_12_2_1),
    .io_keys_12_2_2(dec_io_keys_12_2_2),
    .io_keys_12_2_3(dec_io_keys_12_2_3),
    .io_keys_12_3_0(dec_io_keys_12_3_0),
    .io_keys_12_3_1(dec_io_keys_12_3_1),
    .io_keys_12_3_2(dec_io_keys_12_3_2),
    .io_keys_12_3_3(dec_io_keys_12_3_3),
    .io_keys_13_0_0(dec_io_keys_13_0_0),
    .io_keys_13_0_1(dec_io_keys_13_0_1),
    .io_keys_13_0_2(dec_io_keys_13_0_2),
    .io_keys_13_0_3(dec_io_keys_13_0_3),
    .io_keys_13_1_0(dec_io_keys_13_1_0),
    .io_keys_13_1_1(dec_io_keys_13_1_1),
    .io_keys_13_1_2(dec_io_keys_13_1_2),
    .io_keys_13_1_3(dec_io_keys_13_1_3),
    .io_keys_13_2_0(dec_io_keys_13_2_0),
    .io_keys_13_2_1(dec_io_keys_13_2_1),
    .io_keys_13_2_2(dec_io_keys_13_2_2),
    .io_keys_13_2_3(dec_io_keys_13_2_3),
    .io_keys_13_3_0(dec_io_keys_13_3_0),
    .io_keys_13_3_1(dec_io_keys_13_3_1),
    .io_keys_13_3_2(dec_io_keys_13_3_2),
    .io_keys_13_3_3(dec_io_keys_13_3_3),
    .io_keys_14_0_0(dec_io_keys_14_0_0),
    .io_keys_14_0_1(dec_io_keys_14_0_1),
    .io_keys_14_0_2(dec_io_keys_14_0_2),
    .io_keys_14_0_3(dec_io_keys_14_0_3),
    .io_keys_14_1_0(dec_io_keys_14_1_0),
    .io_keys_14_1_1(dec_io_keys_14_1_1),
    .io_keys_14_1_2(dec_io_keys_14_1_2),
    .io_keys_14_1_3(dec_io_keys_14_1_3),
    .io_keys_14_2_0(dec_io_keys_14_2_0),
    .io_keys_14_2_1(dec_io_keys_14_2_1),
    .io_keys_14_2_2(dec_io_keys_14_2_2),
    .io_keys_14_2_3(dec_io_keys_14_2_3),
    .io_keys_14_3_0(dec_io_keys_14_3_0),
    .io_keys_14_3_1(dec_io_keys_14_3_1),
    .io_keys_14_3_2(dec_io_keys_14_3_2),
    .io_keys_14_3_3(dec_io_keys_14_3_3),
    .io_aes256(dec_io_aes256),
    .io_shiftCyc(dec_io_shiftCyc),
    .io_shiftRev(dec_io_shiftRev),
    .io_shift(dec_io_shift),
    .io_ready(dec_io_ready),
    .io_dataOut(dec_io_dataOut),
    .io_ivOut(dec_io_ivOut),
    .io_outputValid(dec_io_outputValid)
  );
  assign io_encReady = _T_1495 & _T_1496; // @[AesCombined.scala 91:17]
  assign io_decReady = _T_1499 & _T_1496; // @[AesCombined.scala 104:17]
  assign io_encDataOut = enc_io_dataOut; // @[AesCombined.scala 92:19]
  assign io_encIvOut = enc_io_ivOut; // @[AesCombined.scala 93:17]
  assign io_encOutputValid = enc_io_outputValid; // @[AesCombined.scala 94:23]
  assign io_decDataOut = dec_io_dataOut; // @[AesCombined.scala 105:19]
  assign io_decIvOut = dec_io_ivOut; // @[AesCombined.scala 106:17]
  assign io_decOutputValid = dec_io_outputValid; // @[AesCombined.scala 107:23]
  assign shreg_clock = clock;
  assign shreg_io_input = keyUpdate ? _T_1178 : _GEN_3; // @[AesCombined.scala 58:20 AesCombined.scala 68:24 AesCombined.scala 79:24]
  assign shreg_io_enable = _T_1504 | _GEN_39; // @[AesCombined.scala 59:21 AesCombined.scala 67:25 AesCombined.scala 78:25 AesCombined.scala 111:59]
  assign shreg_io_rev = dec_io_shiftRev; // @[AesCombined.scala 110:18]
  assign shreg_io_cyc = enc_io_shiftCyc | dec_io_shiftCyc; // @[AesCombined.scala 109:18]
  assign shreg_io_tap = io_aes256; // @[AesCombined.scala 56:18]
  assign enc_clock = clock;
  assign enc_reset = reset;
  assign enc_io_dataIn = io_encDataIn; // @[AesCombined.scala 85:19]
  assign enc_io_ivIn = io_encIvIn; // @[AesCombined.scala 86:17]
  assign enc_io_dataValid = io_encDataValid; // @[AesCombined.scala 87:22]
  assign enc_io_keys_0_0_0 = shreg_io_output_14[127:120]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_0_1 = shreg_io_output_14[119:112]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_0_2 = shreg_io_output_14[111:104]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_0_3 = shreg_io_output_14[103:96]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_1_0 = shreg_io_output_14[95:88]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_1_1 = shreg_io_output_14[87:80]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_1_2 = shreg_io_output_14[79:72]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_1_3 = shreg_io_output_14[71:64]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_2_0 = shreg_io_output_14[63:56]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_2_1 = shreg_io_output_14[55:48]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_2_2 = shreg_io_output_14[47:40]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_2_3 = shreg_io_output_14[39:32]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_3_0 = shreg_io_output_14[31:24]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_3_1 = shreg_io_output_14[23:16]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_3_2 = shreg_io_output_14[15:8]; // @[AesCombined.scala 88:17]
  assign enc_io_keys_0_3_3 = shreg_io_output_14[7:0]; // @[AesCombined.scala 88:17]
  assign enc_io_aes256 = io_aes256; // @[AesCombined.scala 89:19]
  assign dec_clock = clock;
  assign dec_reset = reset;
  assign dec_io_dataIn = io_decDataIn; // @[AesCombined.scala 98:19]
  assign dec_io_ivIn = io_decIvIn; // @[AesCombined.scala 99:17]
  assign dec_io_dataValid = io_decDataValid; // @[AesCombined.scala 100:22]
  assign dec_io_keys_0_0_0 = shreg_io_output_14[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_0_1 = shreg_io_output_14[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_0_2 = shreg_io_output_14[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_0_3 = shreg_io_output_14[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_1_0 = shreg_io_output_14[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_1_1 = shreg_io_output_14[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_1_2 = shreg_io_output_14[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_1_3 = shreg_io_output_14[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_2_0 = shreg_io_output_14[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_2_1 = shreg_io_output_14[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_2_2 = shreg_io_output_14[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_2_3 = shreg_io_output_14[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_3_0 = shreg_io_output_14[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_3_1 = shreg_io_output_14[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_3_2 = shreg_io_output_14[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_0_3_3 = shreg_io_output_14[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_0_0 = shreg_io_output_13[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_0_1 = shreg_io_output_13[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_0_2 = shreg_io_output_13[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_0_3 = shreg_io_output_13[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_1_0 = shreg_io_output_13[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_1_1 = shreg_io_output_13[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_1_2 = shreg_io_output_13[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_1_3 = shreg_io_output_13[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_2_0 = shreg_io_output_13[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_2_1 = shreg_io_output_13[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_2_2 = shreg_io_output_13[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_2_3 = shreg_io_output_13[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_3_0 = shreg_io_output_13[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_3_1 = shreg_io_output_13[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_3_2 = shreg_io_output_13[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_1_3_3 = shreg_io_output_13[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_0_0 = shreg_io_output_12[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_0_1 = shreg_io_output_12[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_0_2 = shreg_io_output_12[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_0_3 = shreg_io_output_12[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_1_0 = shreg_io_output_12[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_1_1 = shreg_io_output_12[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_1_2 = shreg_io_output_12[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_1_3 = shreg_io_output_12[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_2_0 = shreg_io_output_12[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_2_1 = shreg_io_output_12[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_2_2 = shreg_io_output_12[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_2_3 = shreg_io_output_12[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_3_0 = shreg_io_output_12[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_3_1 = shreg_io_output_12[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_3_2 = shreg_io_output_12[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_2_3_3 = shreg_io_output_12[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_0_0 = shreg_io_output_11[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_0_1 = shreg_io_output_11[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_0_2 = shreg_io_output_11[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_0_3 = shreg_io_output_11[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_1_0 = shreg_io_output_11[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_1_1 = shreg_io_output_11[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_1_2 = shreg_io_output_11[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_1_3 = shreg_io_output_11[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_2_0 = shreg_io_output_11[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_2_1 = shreg_io_output_11[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_2_2 = shreg_io_output_11[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_2_3 = shreg_io_output_11[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_3_0 = shreg_io_output_11[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_3_1 = shreg_io_output_11[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_3_2 = shreg_io_output_11[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_3_3_3 = shreg_io_output_11[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_0_0 = shreg_io_output_10[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_0_1 = shreg_io_output_10[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_0_2 = shreg_io_output_10[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_0_3 = shreg_io_output_10[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_1_0 = shreg_io_output_10[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_1_1 = shreg_io_output_10[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_1_2 = shreg_io_output_10[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_1_3 = shreg_io_output_10[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_2_0 = shreg_io_output_10[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_2_1 = shreg_io_output_10[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_2_2 = shreg_io_output_10[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_2_3 = shreg_io_output_10[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_3_0 = shreg_io_output_10[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_3_1 = shreg_io_output_10[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_3_2 = shreg_io_output_10[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_4_3_3 = shreg_io_output_10[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_0_0 = shreg_io_output_9[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_0_1 = shreg_io_output_9[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_0_2 = shreg_io_output_9[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_0_3 = shreg_io_output_9[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_1_0 = shreg_io_output_9[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_1_1 = shreg_io_output_9[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_1_2 = shreg_io_output_9[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_1_3 = shreg_io_output_9[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_2_0 = shreg_io_output_9[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_2_1 = shreg_io_output_9[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_2_2 = shreg_io_output_9[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_2_3 = shreg_io_output_9[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_3_0 = shreg_io_output_9[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_3_1 = shreg_io_output_9[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_3_2 = shreg_io_output_9[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_5_3_3 = shreg_io_output_9[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_0_0 = shreg_io_output_8[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_0_1 = shreg_io_output_8[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_0_2 = shreg_io_output_8[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_0_3 = shreg_io_output_8[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_1_0 = shreg_io_output_8[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_1_1 = shreg_io_output_8[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_1_2 = shreg_io_output_8[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_1_3 = shreg_io_output_8[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_2_0 = shreg_io_output_8[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_2_1 = shreg_io_output_8[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_2_2 = shreg_io_output_8[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_2_3 = shreg_io_output_8[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_3_0 = shreg_io_output_8[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_3_1 = shreg_io_output_8[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_3_2 = shreg_io_output_8[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_6_3_3 = shreg_io_output_8[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_0_0 = shreg_io_output_7[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_0_1 = shreg_io_output_7[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_0_2 = shreg_io_output_7[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_0_3 = shreg_io_output_7[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_1_0 = shreg_io_output_7[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_1_1 = shreg_io_output_7[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_1_2 = shreg_io_output_7[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_1_3 = shreg_io_output_7[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_2_0 = shreg_io_output_7[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_2_1 = shreg_io_output_7[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_2_2 = shreg_io_output_7[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_2_3 = shreg_io_output_7[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_3_0 = shreg_io_output_7[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_3_1 = shreg_io_output_7[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_3_2 = shreg_io_output_7[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_7_3_3 = shreg_io_output_7[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_0_0 = shreg_io_output_6[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_0_1 = shreg_io_output_6[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_0_2 = shreg_io_output_6[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_0_3 = shreg_io_output_6[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_1_0 = shreg_io_output_6[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_1_1 = shreg_io_output_6[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_1_2 = shreg_io_output_6[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_1_3 = shreg_io_output_6[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_2_0 = shreg_io_output_6[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_2_1 = shreg_io_output_6[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_2_2 = shreg_io_output_6[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_2_3 = shreg_io_output_6[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_3_0 = shreg_io_output_6[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_3_1 = shreg_io_output_6[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_3_2 = shreg_io_output_6[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_8_3_3 = shreg_io_output_6[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_0_0 = shreg_io_output_5[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_0_1 = shreg_io_output_5[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_0_2 = shreg_io_output_5[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_0_3 = shreg_io_output_5[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_1_0 = shreg_io_output_5[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_1_1 = shreg_io_output_5[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_1_2 = shreg_io_output_5[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_1_3 = shreg_io_output_5[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_2_0 = shreg_io_output_5[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_2_1 = shreg_io_output_5[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_2_2 = shreg_io_output_5[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_2_3 = shreg_io_output_5[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_3_0 = shreg_io_output_5[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_3_1 = shreg_io_output_5[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_3_2 = shreg_io_output_5[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_9_3_3 = shreg_io_output_5[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_0_0 = shreg_io_output_4[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_0_1 = shreg_io_output_4[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_0_2 = shreg_io_output_4[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_0_3 = shreg_io_output_4[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_1_0 = shreg_io_output_4[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_1_1 = shreg_io_output_4[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_1_2 = shreg_io_output_4[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_1_3 = shreg_io_output_4[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_2_0 = shreg_io_output_4[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_2_1 = shreg_io_output_4[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_2_2 = shreg_io_output_4[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_2_3 = shreg_io_output_4[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_3_0 = shreg_io_output_4[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_3_1 = shreg_io_output_4[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_3_2 = shreg_io_output_4[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_10_3_3 = shreg_io_output_4[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_0_0 = shreg_io_output_3[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_0_1 = shreg_io_output_3[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_0_2 = shreg_io_output_3[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_0_3 = shreg_io_output_3[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_1_0 = shreg_io_output_3[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_1_1 = shreg_io_output_3[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_1_2 = shreg_io_output_3[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_1_3 = shreg_io_output_3[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_2_0 = shreg_io_output_3[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_2_1 = shreg_io_output_3[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_2_2 = shreg_io_output_3[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_2_3 = shreg_io_output_3[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_3_0 = shreg_io_output_3[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_3_1 = shreg_io_output_3[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_3_2 = shreg_io_output_3[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_11_3_3 = shreg_io_output_3[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_0_0 = shreg_io_output_2[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_0_1 = shreg_io_output_2[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_0_2 = shreg_io_output_2[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_0_3 = shreg_io_output_2[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_1_0 = shreg_io_output_2[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_1_1 = shreg_io_output_2[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_1_2 = shreg_io_output_2[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_1_3 = shreg_io_output_2[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_2_0 = shreg_io_output_2[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_2_1 = shreg_io_output_2[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_2_2 = shreg_io_output_2[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_2_3 = shreg_io_output_2[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_3_0 = shreg_io_output_2[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_3_1 = shreg_io_output_2[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_3_2 = shreg_io_output_2[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_12_3_3 = shreg_io_output_2[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_0_0 = shreg_io_output_1[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_0_1 = shreg_io_output_1[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_0_2 = shreg_io_output_1[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_0_3 = shreg_io_output_1[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_1_0 = shreg_io_output_1[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_1_1 = shreg_io_output_1[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_1_2 = shreg_io_output_1[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_1_3 = shreg_io_output_1[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_2_0 = shreg_io_output_1[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_2_1 = shreg_io_output_1[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_2_2 = shreg_io_output_1[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_2_3 = shreg_io_output_1[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_3_0 = shreg_io_output_1[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_3_1 = shreg_io_output_1[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_3_2 = shreg_io_output_1[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_13_3_3 = shreg_io_output_1[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_0_0 = shreg_io_output_0[127:120]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_0_1 = shreg_io_output_0[119:112]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_0_2 = shreg_io_output_0[111:104]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_0_3 = shreg_io_output_0[103:96]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_1_0 = shreg_io_output_0[95:88]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_1_1 = shreg_io_output_0[87:80]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_1_2 = shreg_io_output_0[79:72]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_1_3 = shreg_io_output_0[71:64]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_2_0 = shreg_io_output_0[63:56]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_2_1 = shreg_io_output_0[55:48]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_2_2 = shreg_io_output_0[47:40]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_2_3 = shreg_io_output_0[39:32]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_3_0 = shreg_io_output_0[31:24]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_3_1 = shreg_io_output_0[23:16]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_3_2 = shreg_io_output_0[15:8]; // @[AesCombined.scala 101:17]
  assign dec_io_keys_14_3_3 = shreg_io_output_0[7:0]; // @[AesCombined.scala 101:17]
  assign dec_io_aes256 = io_aes256; // @[AesCombined.scala 102:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  keyUpdate = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  keyInd = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      keyUpdate <= 1'h0;
    end else if (keyUpdate) begin
      if (_T_6) begin
        keyUpdate <= 1'h0;
      end else begin
        keyUpdate <= _GEN_0;
      end
    end else begin
      keyUpdate <= _GEN_0;
    end
    if (reset) begin
      keyInd <= 6'h0;
    end else if (keyUpdate) begin
      keyInd <= _T_2;
    end else if (io_keyValid) begin
      keyInd <= 6'h1;
    end
  end
endmodule
module AesWishbone(
  input         clock,
  input         reset,
  input         io_bus_cyc,
  input         io_bus_stb,
  input         io_bus_we,
  input  [3:0]  io_bus_sel,
  input  [31:0] io_bus_addr,
  input  [31:0] io_bus_data_wr,
  output        io_bus_ack,
  output [31:0] io_bus_data_rd
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  accel_clock; // @[AesWishbone.scala 38:23]
  wire  accel_reset; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_encDataIn; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_encIvIn; // @[AesWishbone.scala 38:23]
  wire  accel_io_encDataValid; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_decDataIn; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_decIvIn; // @[AesWishbone.scala 38:23]
  wire  accel_io_decDataValid; // @[AesWishbone.scala 38:23]
  wire  accel_io_aes256; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_keyIn; // @[AesWishbone.scala 38:23]
  wire  accel_io_keyShift; // @[AesWishbone.scala 38:23]
  wire  accel_io_keyValid; // @[AesWishbone.scala 38:23]
  wire  accel_io_encReady; // @[AesWishbone.scala 38:23]
  wire  accel_io_decReady; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_encDataOut; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_encIvOut; // @[AesWishbone.scala 38:23]
  wire  accel_io_encOutputValid; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_decDataOut; // @[AesWishbone.scala 38:23]
  wire [127:0] accel_io_decIvOut; // @[AesWishbone.scala 38:23]
  wire  accel_io_decOutputValid; // @[AesWishbone.scala 38:23]
  reg [31:0] data_rd; // @[AesWishbone.scala 31:26]
  reg  ack; // @[AesWishbone.scala 34:22]
  reg  cbcMode; // @[AesWishbone.scala 40:26]
  reg  aes256Mode; // @[AesWishbone.scala 41:29]
  reg [127:0] iv; // @[AesWishbone.scala 42:17]
  reg  outValid; // @[AesWishbone.scala 44:27]
  reg [127:0] out; // @[AesWishbone.scala 45:18]
  reg  _T; // @[RisingEdge.scala 20:45]
  wire  _T_1 = ~_T; // @[RisingEdge.scala 20:37]
  wire  _T_2 = accel_io_encOutputValid & _T_1; // @[RisingEdge.scala 20:34]
  wire  _GEN_1 = _T_2 | outValid; // @[AesWishbone.scala 47:48]
  wire [127:0] _GEN_2 = _T_2 ? accel_io_encIvOut : iv; // @[AesWishbone.scala 47:48]
  reg  _T_3; // @[RisingEdge.scala 20:45]
  wire  _T_4 = ~_T_3; // @[RisingEdge.scala 20:37]
  wire  _T_5 = accel_io_decOutputValid & _T_4; // @[RisingEdge.scala 20:34]
  wire  _GEN_4 = _T_5 | _GEN_1; // @[AesWishbone.scala 53:48]
  wire [127:0] _GEN_5 = _T_5 ? accel_io_decIvOut : _GEN_2; // @[AesWishbone.scala 53:48]
  reg [127:0] dataReg; // @[AesWishbone.scala 59:22]
  wire [31:0] statusReg = {27'h0,aes256Mode,cbcMode,outValid,accel_io_encReady,accel_io_decReady}; // @[Cat.scala 29:58]
  reg [127:0] key; // @[AesWishbone.scala 79:67]
  reg  keyUpdated; // @[AesWishbone.scala 81:29]
  reg  keyShift; // @[AesWishbone.scala 82:27]
  wire  _T_13 = io_bus_cyc & io_bus_stb; // @[AesWishbone.scala 119:21]
  wire  _T_14 = ~io_bus_ack; // @[AesWishbone.scala 119:38]
  wire  _T_15 = _T_13 & _T_14; // @[AesWishbone.scala 119:35]
  wire  _T_35 = 30'h0 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_40 = 30'h1 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_43 = io_bus_sel[0] & io_bus_data_wr[0]; // @[AesWishbone.scala 148:41]
  wire  _T_44 = _T_43 & accel_io_encReady; // @[AesWishbone.scala 148:62]
  wire  _GEN_39 = _T_40 & _T_44; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_35 ? 1'h0 : _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_57 = io_bus_we & _GEN_48; // @[AesWishbone.scala 139:25]
  wire  startEnc = _T_15 & _GEN_57; // @[AesWishbone.scala 119:51]
  wire  _T_45 = 30'h2 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_49 = _T_43 & accel_io_decReady; // @[AesWishbone.scala 152:62]
  wire  _GEN_33 = _T_45 & _T_49; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_40 ? 1'h0 : _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_49 = _T_35 ? 1'h0 : _GEN_40; // @[Conditional.scala 40:58]
  wire  _GEN_58 = io_bus_we & _GEN_49; // @[AesWishbone.scala 139:25]
  wire  startDec = _T_15 & _GEN_58; // @[AesWishbone.scala 119:51]
  wire  _T_12 = startEnc | startDec; // @[AesWishbone.scala 111:20]
  wire  _T_18 = 30'hc == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_20 = 30'hd == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_22 = 30'he == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_24 = 30'hf == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_27 = io_bus_addr[31:2] == 30'h14; // @[AesWishbone.scala 134:44]
  wire  _T_29 = io_bus_addr[31:2] == 30'h15; // @[AesWishbone.scala 134:44]
  wire  _T_31 = io_bus_addr[31:2] == 30'h16; // @[AesWishbone.scala 134:44]
  wire  _T_33 = io_bus_addr[31:2] == 30'h17; // @[AesWishbone.scala 134:44]
  wire  _T_50 = 30'h3 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_55 = _T_49 & accel_io_encReady; // @[AesWishbone.scala 156:74]
  wire  _T_58 = io_bus_sel[0] & io_bus_data_wr[1]; // @[AesWishbone.scala 157:41]
  wire  _T_59 = _T_58 & accel_io_decReady; // @[AesWishbone.scala 157:62]
  wire  _T_60 = _T_59 & accel_io_encReady; // @[AesWishbone.scala 157:74]
  wire  _T_61 = 30'h4 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire [127:0] _T_63 = {dataReg[95:0],io_bus_data_wr}; // @[Cat.scala 29:58]
  wire  _T_64 = 30'h8 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire [127:0] _T_66 = {iv[95:0],io_bus_data_wr}; // @[Cat.scala 29:58]
  wire  _T_67 = 30'h10 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire [127:0] _T_69 = {key[95:0],io_bus_data_wr}; // @[Cat.scala 29:58]
  wire  _GEN_28 = _T_50 & _T_55; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_50 & _T_60; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_45 ? 1'h0 : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_35 = _T_45 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_40 ? 1'h0 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_40 ? 1'h0 : _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_50 = _T_35 ? 1'h0 : _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_51 = _T_35 ? 1'h0 : _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_59 = io_bus_we & _GEN_50; // @[AesWishbone.scala 139:25]
  wire  _GEN_60 = io_bus_we & _GEN_51; // @[AesWishbone.scala 139:25]
  wire  _GEN_70 = _T_15 & _GEN_59; // @[AesWishbone.scala 119:51]
  wire  _GEN_71 = _T_15 & _GEN_60; // @[AesWishbone.scala 119:51]
  AesCombined accel ( // @[AesWishbone.scala 38:23]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_encDataIn(accel_io_encDataIn),
    .io_encIvIn(accel_io_encIvIn),
    .io_encDataValid(accel_io_encDataValid),
    .io_decDataIn(accel_io_decDataIn),
    .io_decIvIn(accel_io_decIvIn),
    .io_decDataValid(accel_io_decDataValid),
    .io_aes256(accel_io_aes256),
    .io_keyIn(accel_io_keyIn),
    .io_keyShift(accel_io_keyShift),
    .io_keyValid(accel_io_keyValid),
    .io_encReady(accel_io_encReady),
    .io_decReady(accel_io_decReady),
    .io_encDataOut(accel_io_encDataOut),
    .io_encIvOut(accel_io_encIvOut),
    .io_encOutputValid(accel_io_encOutputValid),
    .io_decDataOut(accel_io_decDataOut),
    .io_decIvOut(accel_io_decIvOut),
    .io_decOutputValid(accel_io_decOutputValid)
  );
  assign io_bus_ack = ack; // @[AesWishbone.scala 35:16]
  assign io_bus_data_rd = data_rd; // @[AesWishbone.scala 32:20]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_encDataIn = dataReg; // @[AesWishbone.scala 69:24]
  assign accel_io_encIvIn = cbcMode ? iv : 128'h0; // @[AesWishbone.scala 64:22]
  assign accel_io_encDataValid = _T_15 & _GEN_57; // @[AesWishbone.scala 108:27]
  assign accel_io_decDataIn = dataReg; // @[AesWishbone.scala 70:24]
  assign accel_io_decIvIn = cbcMode ? iv : 128'h0; // @[AesWishbone.scala 65:22]
  assign accel_io_decDataValid = _T_15 & _GEN_58; // @[AesWishbone.scala 109:27]
  assign accel_io_aes256 = aes256Mode; // @[AesWishbone.scala 67:21]
  assign accel_io_keyIn = key; // @[AesWishbone.scala 101:20]
  assign accel_io_keyShift = keyShift; // @[AesWishbone.scala 103:23]
  assign accel_io_keyValid = keyUpdated; // @[AesWishbone.scala 102:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_rd = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ack = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cbcMode = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  aes256Mode = _RAND_3[0:0];
  _RAND_4 = {4{`RANDOM}};
  iv = _RAND_4[127:0];
  _RAND_5 = {1{`RANDOM}};
  outValid = _RAND_5[0:0];
  _RAND_6 = {4{`RANDOM}};
  out = _RAND_6[127:0];
  _RAND_7 = {1{`RANDOM}};
  _T = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_3 = _RAND_8[0:0];
  _RAND_9 = {4{`RANDOM}};
  dataReg = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  key = _RAND_10[127:0];
  _RAND_11 = {1{`RANDOM}};
  keyUpdated = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  keyShift = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      data_rd <= 32'h0;
    end else if (_T_15) begin
      if (_T_33) begin
        data_rd <= 32'h65726f;
      end else if (_T_31) begin
        data_rd <= 32'h43203635;
      end else if (_T_29) begin
        data_rd <= 32'h322f3832;
      end else if (_T_27) begin
        data_rd <= 32'h31534541;
      end else if (_T_35) begin
        data_rd <= statusReg;
      end else if (_T_18) begin
        data_rd <= out[127:96];
      end else if (_T_20) begin
        data_rd <= out[95:64];
      end else if (_T_22) begin
        data_rd <= out[63:32];
      end else if (_T_24) begin
        data_rd <= out[31:0];
      end else begin
        data_rd <= 32'h0;
      end
    end
    if (reset) begin
      ack <= 1'h0;
    end else begin
      ack <= _T_15;
    end
    if (reset) begin
      cbcMode <= 1'h0;
    end else if (_T_15) begin
      if (io_bus_we) begin
        if (_T_35) begin
          if (io_bus_sel[0]) begin
            cbcMode <= io_bus_data_wr[3];
          end
        end
      end
    end
    if (reset) begin
      aes256Mode <= 1'h0;
    end else if (_T_15) begin
      if (io_bus_we) begin
        if (_T_35) begin
          if (io_bus_sel[0]) begin
            aes256Mode <= io_bus_data_wr[4];
          end
        end
      end
    end
    if (_T_15) begin
      if (io_bus_we) begin
        if (_T_35) begin
          if (_T_5) begin
            iv <= accel_io_decIvOut;
          end else if (_T_2) begin
            iv <= accel_io_encIvOut;
          end
        end else if (_T_40) begin
          if (_T_5) begin
            iv <= accel_io_decIvOut;
          end else if (_T_2) begin
            iv <= accel_io_encIvOut;
          end
        end else if (_T_45) begin
          if (_T_5) begin
            iv <= accel_io_decIvOut;
          end else if (_T_2) begin
            iv <= accel_io_encIvOut;
          end
        end else if (_T_50) begin
          if (_T_5) begin
            iv <= accel_io_decIvOut;
          end else if (_T_2) begin
            iv <= accel_io_encIvOut;
          end
        end else if (_T_61) begin
          iv <= _GEN_5;
        end else if (_T_64) begin
          iv <= _T_66;
        end else begin
          iv <= _GEN_5;
        end
      end else begin
        iv <= _GEN_5;
      end
    end else begin
      iv <= _GEN_5;
    end
    if (reset) begin
      outValid <= 1'h0;
    end else if (_T_12) begin
      outValid <= 1'h0;
    end else begin
      outValid <= _GEN_4;
    end
    if (_T_5) begin
      out <= accel_io_decDataOut;
    end else if (_T_2) begin
      out <= accel_io_encDataOut;
    end
    _T <= accel_io_encOutputValid;
    _T_3 <= accel_io_decOutputValid;
    if (_T_15) begin
      if (io_bus_we) begin
        if (!(_T_35)) begin
          if (!(_T_40)) begin
            if (!(_T_45)) begin
              if (!(_T_50)) begin
                if (_T_61) begin
                  dataReg <= _T_63;
                end
              end
            end
          end
        end
      end
    end
    if (_T_15) begin
      if (io_bus_we) begin
        if (!(_T_35)) begin
          if (!(_T_40)) begin
            if (!(_T_45)) begin
              if (!(_T_50)) begin
                if (!(_T_61)) begin
                  if (!(_T_64)) begin
                    if (_T_67) begin
                      key <= _T_69;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      keyUpdated <= 1'h0;
    end else begin
      keyUpdated <= _GEN_70;
    end
    if (reset) begin
      keyShift <= 1'h0;
    end else begin
      keyShift <= _GEN_71;
    end
  end
endmodule
module ShiftRegister_1(
  input         clock,
  input  [31:0] io_input,
  input         io_enable,
  output [31:0] io_output_1,
  output [31:0] io_output_6,
  output [31:0] io_output_14,
  output [31:0] io_output_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_0; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_1; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_2; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_3; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_4; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_5; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_6; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_7; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_8; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_9; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_10; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_11; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_12; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_13; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_14; // @[ShiftRegister.scala 34:18]
  reg [31:0] reg_15; // @[ShiftRegister.scala 34:18]
  assign io_output_1 = reg_1; // @[ShiftRegister.scala 53:15]
  assign io_output_6 = reg_6; // @[ShiftRegister.scala 53:15]
  assign io_output_14 = reg_14; // @[ShiftRegister.scala 53:15]
  assign io_output_15 = reg_15; // @[ShiftRegister.scala 53:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_15 = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_enable) begin
      reg_0 <= io_input;
    end
    if (io_enable) begin
      reg_1 <= reg_0;
    end
    if (io_enable) begin
      reg_2 <= reg_1;
    end
    if (io_enable) begin
      reg_3 <= reg_2;
    end
    if (io_enable) begin
      reg_4 <= reg_3;
    end
    if (io_enable) begin
      reg_5 <= reg_4;
    end
    if (io_enable) begin
      reg_6 <= reg_5;
    end
    if (io_enable) begin
      reg_7 <= reg_6;
    end
    if (io_enable) begin
      reg_8 <= reg_7;
    end
    if (io_enable) begin
      reg_9 <= reg_8;
    end
    if (io_enable) begin
      reg_10 <= reg_9;
    end
    if (io_enable) begin
      reg_11 <= reg_10;
    end
    if (io_enable) begin
      reg_12 <= reg_11;
    end
    if (io_enable) begin
      reg_13 <= reg_12;
    end
    if (io_enable) begin
      reg_14 <= reg_13;
    end
    if (io_enable) begin
      reg_15 <= reg_14;
    end
  end
endmodule
module MessageScheduleArray(
  input         clock,
  input         reset,
  input         io_first,
  input         io_shiftIn,
  input  [31:0] io_wordIn,
  output [31:0] io_wOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  shreg_clock; // @[MessageScheduleArray.scala 50:23]
  wire [31:0] shreg_io_input; // @[MessageScheduleArray.scala 50:23]
  wire  shreg_io_enable; // @[MessageScheduleArray.scala 50:23]
  wire [31:0] shreg_io_output_1; // @[MessageScheduleArray.scala 50:23]
  wire [31:0] shreg_io_output_6; // @[MessageScheduleArray.scala 50:23]
  wire [31:0] shreg_io_output_14; // @[MessageScheduleArray.scala 50:23]
  wire [31:0] shreg_io_output_15; // @[MessageScheduleArray.scala 50:23]
  reg [5:0] iReg; // @[MessageScheduleArray.scala 32:23]
  reg [31:0] out; // @[MessageScheduleArray.scala 36:22]
  wire [5:0] _T_1 = iReg + 6'h1; // @[MessageScheduleArray.scala 44:19]
  wire [5:0] _GEN_0 = io_shiftIn ? _T_1 : iReg; // @[MessageScheduleArray.scala 43:30]
  wire [5:0] i = io_first ? 6'h0 : _GEN_0; // @[MessageScheduleArray.scala 40:21]
  wire  _T_4 = i < 6'h10; // @[MessageScheduleArray.scala 60:17]
  wire [31:0] _T_7 = {shreg_io_output_14[6:0],shreg_io_output_14[31:7]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_10 = {shreg_io_output_14[17:0],shreg_io_output_14[31:18]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_11 = _T_7 ^ _T_10; // @[MessageScheduleArray.scala 63:58]
  wire [31:0] _GEN_6 = {{3'd0}, shreg_io_output_14[31:3]}; // @[MessageScheduleArray.scala 63:97]
  wire [31:0] _T_13 = _T_11 ^ _GEN_6; // @[MessageScheduleArray.scala 63:97]
  wire [31:0] _T_16 = {shreg_io_output_1[16:0],shreg_io_output_1[31:17]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_19 = {shreg_io_output_1[18:0],shreg_io_output_1[31:19]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_20 = _T_16 ^ _T_19; // @[MessageScheduleArray.scala 64:58]
  wire [31:0] _GEN_7 = {{10'd0}, shreg_io_output_1[31:10]}; // @[MessageScheduleArray.scala 64:96]
  wire [31:0] _T_22 = _T_20 ^ _GEN_7; // @[MessageScheduleArray.scala 64:96]
  wire [31:0] _T_24 = shreg_io_output_15 + _T_13; // @[MessageScheduleArray.scala 65:44]
  wire [31:0] _T_26 = _T_24 + shreg_io_output_6; // @[MessageScheduleArray.scala 65:49]
  wire [31:0] _T_28 = _T_26 + _T_22; // @[MessageScheduleArray.scala 65:70]
  wire [31:0] _GEN_4 = _T_4 ? io_wordIn : _T_28; // @[MessageScheduleArray.scala 60:25]
  ShiftRegister_1 shreg ( // @[MessageScheduleArray.scala 50:23]
    .clock(shreg_clock),
    .io_input(shreg_io_input),
    .io_enable(shreg_io_enable),
    .io_output_1(shreg_io_output_1),
    .io_output_6(shreg_io_output_6),
    .io_output_14(shreg_io_output_14),
    .io_output_15(shreg_io_output_15)
  );
  assign io_wOut = out; // @[MessageScheduleArray.scala 37:13]
  assign shreg_clock = clock;
  assign shreg_io_input = io_shiftIn ? _GEN_4 : 32'h0; // @[MessageScheduleArray.scala 56:20]
  assign shreg_io_enable = io_shiftIn; // @[MessageScheduleArray.scala 55:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  iReg = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  out = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      iReg <= 6'h0;
    end else if (io_first) begin
      iReg <= 6'h0;
    end else if (io_shiftIn) begin
      iReg <= _T_1;
    end
    if (reset) begin
      out <= 32'h0;
    end else if (io_shiftIn) begin
      if (_T_4) begin
        out <= io_wordIn;
      end else begin
        out <= _T_28;
      end
    end else begin
      out <= 32'h0;
    end
  end
endmodule
module CompressionFunction(
  input         clock,
  input         reset,
  input         io_first,
  input         io_newChunk,
  input         io_shiftIn,
  input  [31:0] io_wordIn,
  output        io_valid,
  output [31:0] io_out_0,
  output [31:0] io_out_1,
  output [31:0] io_out_2,
  output [31:0] io_out_3,
  output [31:0] io_out_4,
  output [31:0] io_out_5,
  output [31:0] io_out_6,
  output [31:0] io_out_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  messageScheduleArray_clock; // @[CompressionFunction.scala 49:38]
  wire  messageScheduleArray_reset; // @[CompressionFunction.scala 49:38]
  wire  messageScheduleArray_io_first; // @[CompressionFunction.scala 49:38]
  wire  messageScheduleArray_io_shiftIn; // @[CompressionFunction.scala 49:38]
  wire [31:0] messageScheduleArray_io_wordIn; // @[CompressionFunction.scala 49:38]
  wire [31:0] messageScheduleArray_io_wOut; // @[CompressionFunction.scala 49:38]
  reg  valid; // @[CompressionFunction.scala 32:24]
  reg [5:0] i; // @[CompressionFunction.scala 35:20]
  reg [31:0] hash_val_0; // @[CompressionFunction.scala 37:27]
  reg [31:0] hash_val_1; // @[CompressionFunction.scala 37:27]
  reg [31:0] hash_val_2; // @[CompressionFunction.scala 37:27]
  reg [31:0] hash_val_3; // @[CompressionFunction.scala 37:27]
  reg [31:0] hash_val_4; // @[CompressionFunction.scala 37:27]
  reg [31:0] hash_val_5; // @[CompressionFunction.scala 37:27]
  reg [31:0] hash_val_6; // @[CompressionFunction.scala 37:27]
  reg [31:0] hash_val_7; // @[CompressionFunction.scala 37:27]
  reg [31:0] a; // @[CompressionFunction.scala 40:20]
  reg [31:0] b; // @[CompressionFunction.scala 41:20]
  reg [31:0] c; // @[CompressionFunction.scala 42:20]
  reg [31:0] d; // @[CompressionFunction.scala 43:20]
  reg [31:0] e; // @[CompressionFunction.scala 44:20]
  reg [31:0] f; // @[CompressionFunction.scala 45:20]
  reg [31:0] g; // @[CompressionFunction.scala 46:20]
  reg [31:0] h; // @[CompressionFunction.scala 47:20]
  wire  _T_9 = io_first | io_newChunk; // @[CompressionFunction.scala 50:47]
  reg  shiftIn; // @[CompressionFunction.scala 57:26]
  wire [31:0] _T_22 = {e[5:0],e[31:6]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_25 = {e[10:0],e[31:11]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_26 = _T_22 ^ _T_25; // @[CompressionFunction.scala 89:36]
  wire [31:0] _T_29 = {e[24:0],e[31:25]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_30 = _T_26 ^ _T_29; // @[CompressionFunction.scala 89:57]
  wire [31:0] _T_31 = e & f; // @[CompressionFunction.scala 90:21]
  wire [31:0] _T_32 = ~e; // @[CompressionFunction.scala 90:30]
  wire [31:0] _T_33 = _T_32 & g; // @[CompressionFunction.scala 90:41]
  wire [31:0] _T_34 = _T_31 ^ _T_33; // @[CompressionFunction.scala 90:26]
  wire [31:0] _T_36 = h + _T_30; // @[CompressionFunction.scala 91:23]
  wire [31:0] _T_38 = _T_36 + _T_34; // @[CompressionFunction.scala 91:28]
  wire [31:0] _GEN_27 = 6'h1 == i ? 32'h71374491 : 32'h428a2f98; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_28 = 6'h2 == i ? 32'hb5c0fbcf : _GEN_27; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_29 = 6'h3 == i ? 32'he9b5dba5 : _GEN_28; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_30 = 6'h4 == i ? 32'h3956c25b : _GEN_29; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_31 = 6'h5 == i ? 32'h59f111f1 : _GEN_30; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_32 = 6'h6 == i ? 32'h923f82a4 : _GEN_31; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_33 = 6'h7 == i ? 32'hab1c5ed5 : _GEN_32; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_34 = 6'h8 == i ? 32'hd807aa98 : _GEN_33; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_35 = 6'h9 == i ? 32'h12835b01 : _GEN_34; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_36 = 6'ha == i ? 32'h243185be : _GEN_35; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_37 = 6'hb == i ? 32'h550c7dc3 : _GEN_36; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_38 = 6'hc == i ? 32'h72be5d74 : _GEN_37; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_39 = 6'hd == i ? 32'h80deb1fe : _GEN_38; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_40 = 6'he == i ? 32'h9bdc06a7 : _GEN_39; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_41 = 6'hf == i ? 32'hc19bf174 : _GEN_40; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_42 = 6'h10 == i ? 32'he49b69c1 : _GEN_41; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_43 = 6'h11 == i ? 32'hefbe4786 : _GEN_42; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_44 = 6'h12 == i ? 32'hfc19dc6 : _GEN_43; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_45 = 6'h13 == i ? 32'h240ca1cc : _GEN_44; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_46 = 6'h14 == i ? 32'h2de92c6f : _GEN_45; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_47 = 6'h15 == i ? 32'h4a7484aa : _GEN_46; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_48 = 6'h16 == i ? 32'h5cb0a9dc : _GEN_47; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_49 = 6'h17 == i ? 32'h76f988da : _GEN_48; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_50 = 6'h18 == i ? 32'h983e5152 : _GEN_49; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_51 = 6'h19 == i ? 32'ha831c66d : _GEN_50; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_52 = 6'h1a == i ? 32'hb00327c8 : _GEN_51; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_53 = 6'h1b == i ? 32'hbf597fc7 : _GEN_52; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_54 = 6'h1c == i ? 32'hc6e00bf3 : _GEN_53; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_55 = 6'h1d == i ? 32'hd5a79147 : _GEN_54; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_56 = 6'h1e == i ? 32'h6ca6351 : _GEN_55; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_57 = 6'h1f == i ? 32'h14292967 : _GEN_56; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_58 = 6'h20 == i ? 32'h27b70a85 : _GEN_57; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_59 = 6'h21 == i ? 32'h2e1b2138 : _GEN_58; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_60 = 6'h22 == i ? 32'h4d2c6dfc : _GEN_59; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_61 = 6'h23 == i ? 32'h53380d13 : _GEN_60; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_62 = 6'h24 == i ? 32'h650a7354 : _GEN_61; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_63 = 6'h25 == i ? 32'h766a0abb : _GEN_62; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_64 = 6'h26 == i ? 32'h81c2c92e : _GEN_63; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_65 = 6'h27 == i ? 32'h92722c85 : _GEN_64; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_66 = 6'h28 == i ? 32'ha2bfe8a1 : _GEN_65; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_67 = 6'h29 == i ? 32'ha81a664b : _GEN_66; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_68 = 6'h2a == i ? 32'hc24b8b70 : _GEN_67; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_69 = 6'h2b == i ? 32'hc76c51a3 : _GEN_68; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_70 = 6'h2c == i ? 32'hd192e819 : _GEN_69; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_71 = 6'h2d == i ? 32'hd6990624 : _GEN_70; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_72 = 6'h2e == i ? 32'hf40e3585 : _GEN_71; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_73 = 6'h2f == i ? 32'h106aa070 : _GEN_72; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_74 = 6'h30 == i ? 32'h19a4c116 : _GEN_73; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_75 = 6'h31 == i ? 32'h1e376c08 : _GEN_74; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_76 = 6'h32 == i ? 32'h2748774c : _GEN_75; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_77 = 6'h33 == i ? 32'h34b0bcb5 : _GEN_76; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_78 = 6'h34 == i ? 32'h391c0cb3 : _GEN_77; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_79 = 6'h35 == i ? 32'h4ed8aa4a : _GEN_78; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_80 = 6'h36 == i ? 32'h5b9cca4f : _GEN_79; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_81 = 6'h37 == i ? 32'h682e6ff3 : _GEN_80; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_82 = 6'h38 == i ? 32'h748f82ee : _GEN_81; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_83 = 6'h39 == i ? 32'h78a5636f : _GEN_82; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_84 = 6'h3a == i ? 32'h84c87814 : _GEN_83; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_85 = 6'h3b == i ? 32'h8cc70208 : _GEN_84; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_86 = 6'h3c == i ? 32'h90befffa : _GEN_85; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_87 = 6'h3d == i ? 32'ha4506ceb : _GEN_86; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_88 = 6'h3e == i ? 32'hbef9a3f7 : _GEN_87; // @[CompressionFunction.scala 91:33]
  wire [31:0] _GEN_89 = 6'h3f == i ? 32'hc67178f2 : _GEN_88; // @[CompressionFunction.scala 91:33]
  wire [31:0] _T_41 = _T_38 + _GEN_89; // @[CompressionFunction.scala 91:33]
  wire [31:0] _T_43 = _T_41 + messageScheduleArray_io_wOut; // @[CompressionFunction.scala 91:69]
  wire [31:0] _T_46 = {a[1:0],a[31:2]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_49 = {a[12:0],a[31:13]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_50 = _T_46 ^ _T_49; // @[CompressionFunction.scala 92:36]
  wire [31:0] _T_53 = {a[21:0],a[31:22]}; // @[RotateLeft.scala 24:38]
  wire [31:0] _T_54 = _T_50 ^ _T_53; // @[CompressionFunction.scala 92:57]
  wire [31:0] _T_55 = a & b; // @[CompressionFunction.scala 93:22]
  wire [31:0] _T_56 = a & c; // @[CompressionFunction.scala 93:32]
  wire [31:0] _T_57 = _T_55 ^ _T_56; // @[CompressionFunction.scala 93:27]
  wire [31:0] _T_58 = b & c; // @[CompressionFunction.scala 93:42]
  wire [31:0] _T_59 = _T_57 ^ _T_58; // @[CompressionFunction.scala 93:37]
  wire [31:0] _T_61 = _T_54 + _T_59; // @[CompressionFunction.scala 94:24]
  wire [31:0] _T_63 = d + _T_43; // @[CompressionFunction.scala 99:16]
  wire [31:0] _T_65 = _T_43 + _T_61; // @[CompressionFunction.scala 103:20]
  wire [5:0] _T_67 = i + 6'h1; // @[CompressionFunction.scala 105:20]
  wire  _T_68 = i == 6'h3f; // @[CompressionFunction.scala 107:17]
  wire [31:0] _T_72 = _T_65 + hash_val_0; // @[CompressionFunction.scala 110:32]
  wire [31:0] _T_74 = a + hash_val_1; // @[CompressionFunction.scala 111:20]
  wire [31:0] _T_76 = b + hash_val_2; // @[CompressionFunction.scala 112:20]
  wire [31:0] _T_78 = c + hash_val_3; // @[CompressionFunction.scala 113:20]
  wire [31:0] _T_82 = _T_63 + hash_val_4; // @[CompressionFunction.scala 114:28]
  wire [31:0] _T_84 = e + hash_val_5; // @[CompressionFunction.scala 115:20]
  wire [31:0] _T_86 = f + hash_val_6; // @[CompressionFunction.scala 116:20]
  wire [31:0] _T_88 = g + hash_val_7; // @[CompressionFunction.scala 117:20]
  wire [31:0] _T_90 = hash_val_0 + _T_43; // @[CompressionFunction.scala 119:40]
  wire [31:0] _T_92 = _T_90 + _T_61; // @[CompressionFunction.scala 119:48]
  wire [31:0] _T_94 = hash_val_1 + a; // @[CompressionFunction.scala 120:40]
  wire [31:0] _T_96 = hash_val_2 + b; // @[CompressionFunction.scala 121:40]
  wire [31:0] _T_98 = hash_val_3 + c; // @[CompressionFunction.scala 122:40]
  wire [31:0] _T_100 = hash_val_4 + d; // @[CompressionFunction.scala 123:40]
  wire [31:0] _T_102 = _T_100 + _T_43; // @[CompressionFunction.scala 123:44]
  wire [31:0] _T_104 = hash_val_5 + e; // @[CompressionFunction.scala 124:40]
  wire [31:0] _T_106 = hash_val_6 + f; // @[CompressionFunction.scala 125:40]
  wire [31:0] _T_108 = hash_val_7 + g; // @[CompressionFunction.scala 126:40]
  MessageScheduleArray messageScheduleArray ( // @[CompressionFunction.scala 49:38]
    .clock(messageScheduleArray_clock),
    .reset(messageScheduleArray_reset),
    .io_first(messageScheduleArray_io_first),
    .io_shiftIn(messageScheduleArray_io_shiftIn),
    .io_wordIn(messageScheduleArray_io_wordIn),
    .io_wOut(messageScheduleArray_io_wOut)
  );
  assign io_valid = valid; // @[CompressionFunction.scala 33:14]
  assign io_out_0 = hash_val_0; // @[CompressionFunction.scala 38:12]
  assign io_out_1 = hash_val_1; // @[CompressionFunction.scala 38:12]
  assign io_out_2 = hash_val_2; // @[CompressionFunction.scala 38:12]
  assign io_out_3 = hash_val_3; // @[CompressionFunction.scala 38:12]
  assign io_out_4 = hash_val_4; // @[CompressionFunction.scala 38:12]
  assign io_out_5 = hash_val_5; // @[CompressionFunction.scala 38:12]
  assign io_out_6 = hash_val_6; // @[CompressionFunction.scala 38:12]
  assign io_out_7 = hash_val_7; // @[CompressionFunction.scala 38:12]
  assign messageScheduleArray_clock = clock;
  assign messageScheduleArray_reset = reset;
  assign messageScheduleArray_io_first = io_first | io_newChunk; // @[CompressionFunction.scala 50:35]
  assign messageScheduleArray_io_shiftIn = io_shiftIn; // @[CompressionFunction.scala 51:37]
  assign messageScheduleArray_io_wordIn = io_wordIn; // @[CompressionFunction.scala 52:36]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  i = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  hash_val_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  hash_val_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  hash_val_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  hash_val_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  hash_val_4 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  hash_val_5 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  hash_val_6 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hash_val_7 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  a = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  b = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  c = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  d = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  e = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  f = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  g = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  h = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  shiftIn = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      valid <= 1'h0;
    end else if (shiftIn) begin
      valid <= _T_68;
    end else if (_T_9) begin
      valid <= 1'h0;
    end
    if (reset) begin
      i <= 6'h0;
    end else if (shiftIn) begin
      i <= _T_67;
    end else if (_T_9) begin
      i <= 6'h0;
    end
    if (reset) begin
      hash_val_0 <= 32'h6a09e667;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_0 <= _T_92;
      end else if (io_first) begin
        hash_val_0 <= 32'h6a09e667;
      end
    end else if (io_first) begin
      hash_val_0 <= 32'h6a09e667;
    end
    if (reset) begin
      hash_val_1 <= 32'hbb67ae85;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_1 <= _T_94;
      end else if (io_first) begin
        hash_val_1 <= 32'hbb67ae85;
      end
    end else if (io_first) begin
      hash_val_1 <= 32'hbb67ae85;
    end
    if (reset) begin
      hash_val_2 <= 32'h3c6ef372;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_2 <= _T_96;
      end else if (io_first) begin
        hash_val_2 <= 32'h3c6ef372;
      end
    end else if (io_first) begin
      hash_val_2 <= 32'h3c6ef372;
    end
    if (reset) begin
      hash_val_3 <= 32'ha54ff53a;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_3 <= _T_98;
      end else if (io_first) begin
        hash_val_3 <= 32'ha54ff53a;
      end
    end else if (io_first) begin
      hash_val_3 <= 32'ha54ff53a;
    end
    if (reset) begin
      hash_val_4 <= 32'h510e527f;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_4 <= _T_102;
      end else if (io_first) begin
        hash_val_4 <= 32'h510e527f;
      end
    end else if (io_first) begin
      hash_val_4 <= 32'h510e527f;
    end
    if (reset) begin
      hash_val_5 <= 32'h9b05688c;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_5 <= _T_104;
      end else if (io_first) begin
        hash_val_5 <= 32'h9b05688c;
      end
    end else if (io_first) begin
      hash_val_5 <= 32'h9b05688c;
    end
    if (reset) begin
      hash_val_6 <= 32'h1f83d9ab;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_6 <= _T_106;
      end else if (io_first) begin
        hash_val_6 <= 32'h1f83d9ab;
      end
    end else if (io_first) begin
      hash_val_6 <= 32'h1f83d9ab;
    end
    if (reset) begin
      hash_val_7 <= 32'h5be0cd19;
    end else if (shiftIn) begin
      if (_T_68) begin
        hash_val_7 <= _T_108;
      end else if (io_first) begin
        hash_val_7 <= 32'h5be0cd19;
      end
    end else if (io_first) begin
      hash_val_7 <= 32'h5be0cd19;
    end
    if (reset) begin
      a <= 32'h6a09e667;
    end else if (shiftIn) begin
      if (_T_68) begin
        a <= _T_72;
      end else begin
        a <= _T_65;
      end
    end else if (io_first) begin
      a <= 32'h6a09e667;
    end else if (io_newChunk) begin
      a <= hash_val_0;
    end
    if (reset) begin
      b <= 32'hbb67ae85;
    end else if (shiftIn) begin
      if (_T_68) begin
        b <= _T_74;
      end else begin
        b <= a;
      end
    end else if (io_first) begin
      b <= 32'hbb67ae85;
    end else if (io_newChunk) begin
      b <= hash_val_1;
    end
    if (reset) begin
      c <= 32'h3c6ef372;
    end else if (shiftIn) begin
      if (_T_68) begin
        c <= _T_76;
      end else begin
        c <= b;
      end
    end else if (io_first) begin
      c <= 32'h3c6ef372;
    end else if (io_newChunk) begin
      c <= hash_val_2;
    end
    if (reset) begin
      d <= 32'ha54ff53a;
    end else if (shiftIn) begin
      if (_T_68) begin
        d <= _T_78;
      end else begin
        d <= c;
      end
    end else if (io_first) begin
      d <= 32'ha54ff53a;
    end else if (io_newChunk) begin
      d <= hash_val_3;
    end
    if (reset) begin
      e <= 32'h510e527f;
    end else if (shiftIn) begin
      if (_T_68) begin
        e <= _T_82;
      end else begin
        e <= _T_63;
      end
    end else if (io_first) begin
      e <= 32'h510e527f;
    end else if (io_newChunk) begin
      e <= hash_val_4;
    end
    if (reset) begin
      f <= 32'h9b05688c;
    end else if (shiftIn) begin
      if (_T_68) begin
        f <= _T_84;
      end else begin
        f <= e;
      end
    end else if (io_first) begin
      f <= 32'h9b05688c;
    end else if (io_newChunk) begin
      f <= hash_val_5;
    end
    if (reset) begin
      g <= 32'h1f83d9ab;
    end else if (shiftIn) begin
      if (_T_68) begin
        g <= _T_86;
      end else begin
        g <= f;
      end
    end else if (io_first) begin
      g <= 32'h1f83d9ab;
    end else if (io_newChunk) begin
      g <= hash_val_6;
    end
    if (reset) begin
      h <= 32'h5be0cd19;
    end else if (shiftIn) begin
      if (_T_68) begin
        h <= _T_88;
      end else begin
        h <= g;
      end
    end else if (io_first) begin
      h <= 32'h5be0cd19;
    end else if (io_newChunk) begin
      h <= hash_val_7;
    end
    shiftIn <= io_shiftIn;
  end
endmodule
module Sha256Accel(
  input         clock,
  input         reset,
  input         io_first,
  input  [31:0] io_inputData,
  input         io_inputValid,
  output        io_inputReady,
  output [31:0] io_outputData_0,
  output [31:0] io_outputData_1,
  output [31:0] io_outputData_2,
  output [31:0] io_outputData_3,
  output [31:0] io_outputData_4,
  output [31:0] io_outputData_5,
  output [31:0] io_outputData_6,
  output [31:0] io_outputData_7,
  output        io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  accel_clock; // @[Sha256Accel.scala 35:23]
  wire  accel_reset; // @[Sha256Accel.scala 35:23]
  wire  accel_io_first; // @[Sha256Accel.scala 35:23]
  wire  accel_io_newChunk; // @[Sha256Accel.scala 35:23]
  wire  accel_io_shiftIn; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_wordIn; // @[Sha256Accel.scala 35:23]
  wire  accel_io_valid; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_0; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_1; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_2; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_3; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_4; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_5; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_6; // @[Sha256Accel.scala 35:23]
  wire [31:0] accel_io_out_7; // @[Sha256Accel.scala 35:23]
  reg  first; // @[Sha256Accel.scala 39:24]
  wire  _GEN_0 = io_first | first; // @[Sha256Accel.scala 40:21]
  wire  _GEN_1 = accel_io_shiftIn ? 1'h0 : _GEN_0; // @[Sha256Accel.scala 41:29]
  reg [7:0] ctr; // @[Sha256Accel.scala 43:22]
  wire  _T = ctr == 8'h0; // @[Sha256Accel.scala 44:31]
  reg [7:0] _T_3; // @[Sha256Accel.scala 49:30]
  wire  _T_4 = _T_3 < 8'h10; // @[Sha256Accel.scala 49:36]
  wire  _T_5 = ctr < 8'h10; // @[Sha256Accel.scala 49:52]
  wire  _T_6 = _T_4 & _T_5; // @[Sha256Accel.scala 49:44]
  wire  _T_7 = ~io_first; // @[Sha256Accel.scala 49:63]
  wire  _T_8 = _T_6 & _T_7; // @[Sha256Accel.scala 49:60]
  wire  _T_9 = ctr >= 8'h10; // @[Sha256Accel.scala 50:15]
  wire [7:0] _T_11 = ctr + 8'h1; // @[Sha256Accel.scala 54:20]
  wire  _T_12 = ctr == 8'h3f; // @[Sha256Accel.scala 55:19]
  CompressionFunction accel ( // @[Sha256Accel.scala 35:23]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_first(accel_io_first),
    .io_newChunk(accel_io_newChunk),
    .io_shiftIn(accel_io_shiftIn),
    .io_wordIn(accel_io_wordIn),
    .io_valid(accel_io_valid),
    .io_out_0(accel_io_out_0),
    .io_out_1(accel_io_out_1),
    .io_out_2(accel_io_out_2),
    .io_out_3(accel_io_out_3),
    .io_out_4(accel_io_out_4),
    .io_out_5(accel_io_out_5),
    .io_out_6(accel_io_out_6),
    .io_out_7(accel_io_out_7)
  );
  assign io_inputReady = _T_9 ? 1'h0 : _T_8; // @[Sha256Accel.scala 49:19 Sha256Accel.scala 51:23]
  assign io_outputData_0 = accel_io_out_0; // @[Sha256Accel.scala 36:19]
  assign io_outputData_1 = accel_io_out_1; // @[Sha256Accel.scala 36:19]
  assign io_outputData_2 = accel_io_out_2; // @[Sha256Accel.scala 36:19]
  assign io_outputData_3 = accel_io_out_3; // @[Sha256Accel.scala 36:19]
  assign io_outputData_4 = accel_io_out_4; // @[Sha256Accel.scala 36:19]
  assign io_outputData_5 = accel_io_out_5; // @[Sha256Accel.scala 36:19]
  assign io_outputData_6 = accel_io_out_6; // @[Sha256Accel.scala 36:19]
  assign io_outputData_7 = accel_io_out_7; // @[Sha256Accel.scala 36:19]
  assign io_outputValid = accel_io_valid; // @[Sha256Accel.scala 37:20]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_first = first & accel_io_shiftIn; // @[Sha256Accel.scala 45:20]
  assign accel_io_newChunk = _T & accel_io_shiftIn; // @[Sha256Accel.scala 44:23]
  assign accel_io_shiftIn = _T_9 | io_inputValid; // @[Sha256Accel.scala 47:22 Sha256Accel.scala 52:26 Sha256Accel.scala 57:26]
  assign accel_io_wordIn = io_inputData; // @[Sha256Accel.scala 48:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  first = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ctr = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    first <= reset | _GEN_1;
    if (reset) begin
      ctr <= 8'h0;
    end else if (io_first) begin
      ctr <= 8'h0;
    end else if (_T_9) begin
      if (_T_12) begin
        ctr <= 8'h0;
      end else begin
        ctr <= _T_11;
      end
    end else if (io_inputValid) begin
      ctr <= _T_11;
    end
    _T_3 <= ctr;
  end
endmodule
module Sha256Wishbone(
  input         clock,
  input         reset,
  input         io_bus_cyc,
  input         io_bus_stb,
  input         io_bus_we,
  input  [3:0]  io_bus_sel,
  input  [31:0] io_bus_addr,
  input  [31:0] io_bus_data_wr,
  output        io_bus_ack,
  output [31:0] io_bus_data_rd
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  accel_clock; // @[Sha256Wishbone.scala 54:23]
  wire  accel_reset; // @[Sha256Wishbone.scala 54:23]
  wire  accel_io_first; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_inputData; // @[Sha256Wishbone.scala 54:23]
  wire  accel_io_inputValid; // @[Sha256Wishbone.scala 54:23]
  wire  accel_io_inputReady; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_0; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_1; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_2; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_3; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_4; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_5; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_6; // @[Sha256Wishbone.scala 54:23]
  wire [31:0] accel_io_outputData_7; // @[Sha256Wishbone.scala 54:23]
  wire  accel_io_outputValid; // @[Sha256Wishbone.scala 54:23]
  reg [31:0] data_rd; // @[Sha256Wishbone.scala 47:22]
  reg  ack; // @[Sha256Wishbone.scala 50:22]
  wire  _T = io_bus_cyc & io_bus_stb; // @[Sha256Wishbone.scala 61:21]
  wire  _T_1 = ~io_bus_ack; // @[Sha256Wishbone.scala 61:38]
  wire  _T_2 = _T & _T_1; // @[Sha256Wishbone.scala 61:35]
  wire  _T_4 = 30'h0 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_5 = accel_io_outputValid; // @[Sha256Wishbone.scala 65:70]
  wire  _T_6 = accel_io_inputReady; // @[Sha256Wishbone.scala 65:94]
  wire [31:0] _T_9 = {29'h0,_T_5,_T_6,1'h0}; // @[Cat.scala 29:58]
  wire  _T_10 = 30'h4 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_13 = 30'h5 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_16 = 30'h6 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_19 = 30'h7 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_22 = 30'h8 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_25 = 30'h9 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_28 = 30'ha == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_31 = 30'hb == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _T_35 = io_bus_addr[31:2] == 30'h14; // @[Sha256Wishbone.scala 80:44]
  wire  _T_37 = io_bus_addr[31:2] == 30'h15; // @[Sha256Wishbone.scala 80:44]
  wire  _T_39 = io_bus_addr[31:2] == 30'h16; // @[Sha256Wishbone.scala 80:44]
  wire  _T_44 = io_bus_sel[0] & io_bus_data_wr[0]; // @[Sha256Wishbone.scala 90:41]
  wire  _T_45 = 30'h1 == io_bus_addr[31:2]; // @[Conditional.scala 37:30]
  wire  _GEN_14 = _T_45 & _T_6; // @[Conditional.scala 39:67]
  wire  _GEN_15 = _T_45 ? _T_6 : 1'h1; // @[Conditional.scala 39:67]
  wire  _GEN_16 = _T_4 & _T_44; // @[Conditional.scala 40:58]
  wire  _GEN_17 = _T_4 ? 1'h0 : _GEN_14; // @[Conditional.scala 40:58]
  wire  _GEN_18 = _T_4 | _GEN_15; // @[Conditional.scala 40:58]
  wire  _GEN_19 = io_bus_we & _GEN_16; // @[Sha256Wishbone.scala 86:25]
  wire  _GEN_20 = io_bus_we & _GEN_17; // @[Sha256Wishbone.scala 86:25]
  wire  _GEN_21 = io_bus_we ? _GEN_18 : 1'h1; // @[Sha256Wishbone.scala 86:25]
  wire  _GEN_23 = _T_2 & _GEN_21; // @[Sha256Wishbone.scala 61:51]
  Sha256Accel accel ( // @[Sha256Wishbone.scala 54:23]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_first(accel_io_first),
    .io_inputData(accel_io_inputData),
    .io_inputValid(accel_io_inputValid),
    .io_inputReady(accel_io_inputReady),
    .io_outputData_0(accel_io_outputData_0),
    .io_outputData_1(accel_io_outputData_1),
    .io_outputData_2(accel_io_outputData_2),
    .io_outputData_3(accel_io_outputData_3),
    .io_outputData_4(accel_io_outputData_4),
    .io_outputData_5(accel_io_outputData_5),
    .io_outputData_6(accel_io_outputData_6),
    .io_outputData_7(accel_io_outputData_7),
    .io_outputValid(accel_io_outputValid)
  );
  assign io_bus_ack = ack; // @[Sha256Wishbone.scala 51:16]
  assign io_bus_data_rd = data_rd; // @[Sha256Wishbone.scala 48:20]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_first = _T_2 & _GEN_19; // @[Sha256Wishbone.scala 58:20 Sha256Wishbone.scala 91:40]
  assign accel_io_inputData = io_bus_data_wr; // @[Sha256Wishbone.scala 57:24]
  assign accel_io_inputValid = _T_2 & _GEN_20; // @[Sha256Wishbone.scala 56:25 Sha256Wishbone.scala 98:45]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_rd = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ack = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_2) begin
      if (_T_39) begin
        data_rd <= 32'h65726f;
      end else if (_T_37) begin
        data_rd <= 32'h43203635;
      end else if (_T_35) begin
        data_rd <= 32'h32414853;
      end else if (_T_4) begin
        data_rd <= _T_9;
      end else if (_T_10) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_0;
        end else begin
          data_rd <= 32'h0;
        end
      end else if (_T_13) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_1;
        end else begin
          data_rd <= 32'h0;
        end
      end else if (_T_16) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_2;
        end else begin
          data_rd <= 32'h0;
        end
      end else if (_T_19) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_3;
        end else begin
          data_rd <= 32'h0;
        end
      end else if (_T_22) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_4;
        end else begin
          data_rd <= 32'h0;
        end
      end else if (_T_25) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_5;
        end else begin
          data_rd <= 32'h0;
        end
      end else if (_T_28) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_6;
        end else begin
          data_rd <= 32'h0;
        end
      end else if (_T_31) begin
        if (_T_5) begin
          data_rd <= accel_io_outputData_7;
        end else begin
          data_rd <= 32'h0;
        end
      end else begin
        data_rd <= 32'h0;
      end
    end
    if (reset) begin
      ack <= 1'h0;
    end else begin
      ack <= _GEN_23;
    end
  end
endmodule
module AcceleratorTop(
  input         clock,
  input         reset,
  input         io_bus_cyc,
  input         io_bus_stb,
  input         io_bus_we,
  input  [3:0]  io_bus_sel,
  input  [31:0] io_bus_addr,
  input  [31:0] io_bus_data_wr,
  output        io_bus_ack,
  output        io_bus_err,
  output [31:0] io_bus_data_rd
);
  wire  aes_clock; // @[AcceleratorTop.scala 34:21]
  wire  aes_reset; // @[AcceleratorTop.scala 34:21]
  wire  aes_io_bus_cyc; // @[AcceleratorTop.scala 34:21]
  wire  aes_io_bus_stb; // @[AcceleratorTop.scala 34:21]
  wire  aes_io_bus_we; // @[AcceleratorTop.scala 34:21]
  wire [3:0] aes_io_bus_sel; // @[AcceleratorTop.scala 34:21]
  wire [31:0] aes_io_bus_addr; // @[AcceleratorTop.scala 34:21]
  wire [31:0] aes_io_bus_data_wr; // @[AcceleratorTop.scala 34:21]
  wire  aes_io_bus_ack; // @[AcceleratorTop.scala 34:21]
  wire [31:0] aes_io_bus_data_rd; // @[AcceleratorTop.scala 34:21]
  wire  sha256_clock; // @[AcceleratorTop.scala 43:24]
  wire  sha256_reset; // @[AcceleratorTop.scala 43:24]
  wire  sha256_io_bus_cyc; // @[AcceleratorTop.scala 43:24]
  wire  sha256_io_bus_stb; // @[AcceleratorTop.scala 43:24]
  wire  sha256_io_bus_we; // @[AcceleratorTop.scala 43:24]
  wire [3:0] sha256_io_bus_sel; // @[AcceleratorTop.scala 43:24]
  wire [31:0] sha256_io_bus_addr; // @[AcceleratorTop.scala 43:24]
  wire [31:0] sha256_io_bus_data_wr; // @[AcceleratorTop.scala 43:24]
  wire  sha256_io_bus_ack; // @[AcceleratorTop.scala 43:24]
  wire [31:0] sha256_io_bus_data_rd; // @[AcceleratorTop.scala 43:24]
  wire  _T_2 = io_bus_addr[19:16] == 4'h0; // @[AcceleratorTop.scala 41:58]
  wire  _T_6 = io_bus_addr[19:16] == 4'h1; // @[AcceleratorTop.scala 50:61]
  AesWishbone aes ( // @[AcceleratorTop.scala 34:21]
    .clock(aes_clock),
    .reset(aes_reset),
    .io_bus_cyc(aes_io_bus_cyc),
    .io_bus_stb(aes_io_bus_stb),
    .io_bus_we(aes_io_bus_we),
    .io_bus_sel(aes_io_bus_sel),
    .io_bus_addr(aes_io_bus_addr),
    .io_bus_data_wr(aes_io_bus_data_wr),
    .io_bus_ack(aes_io_bus_ack),
    .io_bus_data_rd(aes_io_bus_data_rd)
  );
  Sha256Wishbone sha256 ( // @[AcceleratorTop.scala 43:24]
    .clock(sha256_clock),
    .reset(sha256_reset),
    .io_bus_cyc(sha256_io_bus_cyc),
    .io_bus_stb(sha256_io_bus_stb),
    .io_bus_we(sha256_io_bus_we),
    .io_bus_sel(sha256_io_bus_sel),
    .io_bus_addr(sha256_io_bus_addr),
    .io_bus_data_wr(sha256_io_bus_data_wr),
    .io_bus_ack(sha256_io_bus_ack),
    .io_bus_data_rd(sha256_io_bus_data_rd)
  );
  assign io_bus_ack = _T_2 ? aes_io_bus_ack : sha256_io_bus_ack; // @[AcceleratorTop.scala 53:16]
  assign io_bus_err = 1'h0; // @[AcceleratorTop.scala 54:16]
  assign io_bus_data_rd = _T_2 ? aes_io_bus_data_rd : sha256_io_bus_data_rd; // @[AcceleratorTop.scala 52:20]
  assign aes_clock = clock;
  assign aes_reset = reset;
  assign aes_io_bus_cyc = io_bus_cyc & _T_2; // @[AcceleratorTop.scala 41:20]
  assign aes_io_bus_stb = io_bus_stb; // @[AcceleratorTop.scala 35:20]
  assign aes_io_bus_we = io_bus_we; // @[AcceleratorTop.scala 36:19]
  assign aes_io_bus_sel = io_bus_sel; // @[AcceleratorTop.scala 37:20]
  assign aes_io_bus_addr = {{16'd0}, io_bus_addr[15:0]}; // @[AcceleratorTop.scala 38:21]
  assign aes_io_bus_data_wr = io_bus_data_wr; // @[AcceleratorTop.scala 39:24]
  assign sha256_clock = clock;
  assign sha256_reset = reset;
  assign sha256_io_bus_cyc = io_bus_cyc & _T_6; // @[AcceleratorTop.scala 50:23]
  assign sha256_io_bus_stb = io_bus_stb; // @[AcceleratorTop.scala 44:23]
  assign sha256_io_bus_we = io_bus_we; // @[AcceleratorTop.scala 45:22]
  assign sha256_io_bus_sel = io_bus_sel; // @[AcceleratorTop.scala 46:23]
  assign sha256_io_bus_addr = {{16'd0}, io_bus_addr[15:0]}; // @[AcceleratorTop.scala 47:24]
  assign sha256_io_bus_data_wr = io_bus_data_wr; // @[AcceleratorTop.scala 48:27]
endmodule
