module CLZ(
  input  [107:0] io_in,
  output [6:0]   io_out
);
  wire [6:0] _T_108 = io_in[1] ? 7'h6a : 7'h6b; // @[Mux.scala 47:69]
  wire [6:0] _T_109 = io_in[2] ? 7'h69 : _T_108; // @[Mux.scala 47:69]
  wire [6:0] _T_110 = io_in[3] ? 7'h68 : _T_109; // @[Mux.scala 47:69]
  wire [6:0] _T_111 = io_in[4] ? 7'h67 : _T_110; // @[Mux.scala 47:69]
  wire [6:0] _T_112 = io_in[5] ? 7'h66 : _T_111; // @[Mux.scala 47:69]
  wire [6:0] _T_113 = io_in[6] ? 7'h65 : _T_112; // @[Mux.scala 47:69]
  wire [6:0] _T_114 = io_in[7] ? 7'h64 : _T_113; // @[Mux.scala 47:69]
  wire [6:0] _T_115 = io_in[8] ? 7'h63 : _T_114; // @[Mux.scala 47:69]
  wire [6:0] _T_116 = io_in[9] ? 7'h62 : _T_115; // @[Mux.scala 47:69]
  wire [6:0] _T_117 = io_in[10] ? 7'h61 : _T_116; // @[Mux.scala 47:69]
  wire [6:0] _T_118 = io_in[11] ? 7'h60 : _T_117; // @[Mux.scala 47:69]
  wire [6:0] _T_119 = io_in[12] ? 7'h5f : _T_118; // @[Mux.scala 47:69]
  wire [6:0] _T_120 = io_in[13] ? 7'h5e : _T_119; // @[Mux.scala 47:69]
  wire [6:0] _T_121 = io_in[14] ? 7'h5d : _T_120; // @[Mux.scala 47:69]
  wire [6:0] _T_122 = io_in[15] ? 7'h5c : _T_121; // @[Mux.scala 47:69]
  wire [6:0] _T_123 = io_in[16] ? 7'h5b : _T_122; // @[Mux.scala 47:69]
  wire [6:0] _T_124 = io_in[17] ? 7'h5a : _T_123; // @[Mux.scala 47:69]
  wire [6:0] _T_125 = io_in[18] ? 7'h59 : _T_124; // @[Mux.scala 47:69]
  wire [6:0] _T_126 = io_in[19] ? 7'h58 : _T_125; // @[Mux.scala 47:69]
  wire [6:0] _T_127 = io_in[20] ? 7'h57 : _T_126; // @[Mux.scala 47:69]
  wire [6:0] _T_128 = io_in[21] ? 7'h56 : _T_127; // @[Mux.scala 47:69]
  wire [6:0] _T_129 = io_in[22] ? 7'h55 : _T_128; // @[Mux.scala 47:69]
  wire [6:0] _T_130 = io_in[23] ? 7'h54 : _T_129; // @[Mux.scala 47:69]
  wire [6:0] _T_131 = io_in[24] ? 7'h53 : _T_130; // @[Mux.scala 47:69]
  wire [6:0] _T_132 = io_in[25] ? 7'h52 : _T_131; // @[Mux.scala 47:69]
  wire [6:0] _T_133 = io_in[26] ? 7'h51 : _T_132; // @[Mux.scala 47:69]
  wire [6:0] _T_134 = io_in[27] ? 7'h50 : _T_133; // @[Mux.scala 47:69]
  wire [6:0] _T_135 = io_in[28] ? 7'h4f : _T_134; // @[Mux.scala 47:69]
  wire [6:0] _T_136 = io_in[29] ? 7'h4e : _T_135; // @[Mux.scala 47:69]
  wire [6:0] _T_137 = io_in[30] ? 7'h4d : _T_136; // @[Mux.scala 47:69]
  wire [6:0] _T_138 = io_in[31] ? 7'h4c : _T_137; // @[Mux.scala 47:69]
  wire [6:0] _T_139 = io_in[32] ? 7'h4b : _T_138; // @[Mux.scala 47:69]
  wire [6:0] _T_140 = io_in[33] ? 7'h4a : _T_139; // @[Mux.scala 47:69]
  wire [6:0] _T_141 = io_in[34] ? 7'h49 : _T_140; // @[Mux.scala 47:69]
  wire [6:0] _T_142 = io_in[35] ? 7'h48 : _T_141; // @[Mux.scala 47:69]
  wire [6:0] _T_143 = io_in[36] ? 7'h47 : _T_142; // @[Mux.scala 47:69]
  wire [6:0] _T_144 = io_in[37] ? 7'h46 : _T_143; // @[Mux.scala 47:69]
  wire [6:0] _T_145 = io_in[38] ? 7'h45 : _T_144; // @[Mux.scala 47:69]
  wire [6:0] _T_146 = io_in[39] ? 7'h44 : _T_145; // @[Mux.scala 47:69]
  wire [6:0] _T_147 = io_in[40] ? 7'h43 : _T_146; // @[Mux.scala 47:69]
  wire [6:0] _T_148 = io_in[41] ? 7'h42 : _T_147; // @[Mux.scala 47:69]
  wire [6:0] _T_149 = io_in[42] ? 7'h41 : _T_148; // @[Mux.scala 47:69]
  wire [6:0] _T_150 = io_in[43] ? 7'h40 : _T_149; // @[Mux.scala 47:69]
  wire [6:0] _T_151 = io_in[44] ? 7'h3f : _T_150; // @[Mux.scala 47:69]
  wire [6:0] _T_152 = io_in[45] ? 7'h3e : _T_151; // @[Mux.scala 47:69]
  wire [6:0] _T_153 = io_in[46] ? 7'h3d : _T_152; // @[Mux.scala 47:69]
  wire [6:0] _T_154 = io_in[47] ? 7'h3c : _T_153; // @[Mux.scala 47:69]
  wire [6:0] _T_155 = io_in[48] ? 7'h3b : _T_154; // @[Mux.scala 47:69]
  wire [6:0] _T_156 = io_in[49] ? 7'h3a : _T_155; // @[Mux.scala 47:69]
  wire [6:0] _T_157 = io_in[50] ? 7'h39 : _T_156; // @[Mux.scala 47:69]
  wire [6:0] _T_158 = io_in[51] ? 7'h38 : _T_157; // @[Mux.scala 47:69]
  wire [6:0] _T_159 = io_in[52] ? 7'h37 : _T_158; // @[Mux.scala 47:69]
  wire [6:0] _T_160 = io_in[53] ? 7'h36 : _T_159; // @[Mux.scala 47:69]
  wire [6:0] _T_161 = io_in[54] ? 7'h35 : _T_160; // @[Mux.scala 47:69]
  wire [6:0] _T_162 = io_in[55] ? 7'h34 : _T_161; // @[Mux.scala 47:69]
  wire [6:0] _T_163 = io_in[56] ? 7'h33 : _T_162; // @[Mux.scala 47:69]
  wire [6:0] _T_164 = io_in[57] ? 7'h32 : _T_163; // @[Mux.scala 47:69]
  wire [6:0] _T_165 = io_in[58] ? 7'h31 : _T_164; // @[Mux.scala 47:69]
  wire [6:0] _T_166 = io_in[59] ? 7'h30 : _T_165; // @[Mux.scala 47:69]
  wire [6:0] _T_167 = io_in[60] ? 7'h2f : _T_166; // @[Mux.scala 47:69]
  wire [6:0] _T_168 = io_in[61] ? 7'h2e : _T_167; // @[Mux.scala 47:69]
  wire [6:0] _T_169 = io_in[62] ? 7'h2d : _T_168; // @[Mux.scala 47:69]
  wire [6:0] _T_170 = io_in[63] ? 7'h2c : _T_169; // @[Mux.scala 47:69]
  wire [6:0] _T_171 = io_in[64] ? 7'h2b : _T_170; // @[Mux.scala 47:69]
  wire [6:0] _T_172 = io_in[65] ? 7'h2a : _T_171; // @[Mux.scala 47:69]
  wire [6:0] _T_173 = io_in[66] ? 7'h29 : _T_172; // @[Mux.scala 47:69]
  wire [6:0] _T_174 = io_in[67] ? 7'h28 : _T_173; // @[Mux.scala 47:69]
  wire [6:0] _T_175 = io_in[68] ? 7'h27 : _T_174; // @[Mux.scala 47:69]
  wire [6:0] _T_176 = io_in[69] ? 7'h26 : _T_175; // @[Mux.scala 47:69]
  wire [6:0] _T_177 = io_in[70] ? 7'h25 : _T_176; // @[Mux.scala 47:69]
  wire [6:0] _T_178 = io_in[71] ? 7'h24 : _T_177; // @[Mux.scala 47:69]
  wire [6:0] _T_179 = io_in[72] ? 7'h23 : _T_178; // @[Mux.scala 47:69]
  wire [6:0] _T_180 = io_in[73] ? 7'h22 : _T_179; // @[Mux.scala 47:69]
  wire [6:0] _T_181 = io_in[74] ? 7'h21 : _T_180; // @[Mux.scala 47:69]
  wire [6:0] _T_182 = io_in[75] ? 7'h20 : _T_181; // @[Mux.scala 47:69]
  wire [6:0] _T_183 = io_in[76] ? 7'h1f : _T_182; // @[Mux.scala 47:69]
  wire [6:0] _T_184 = io_in[77] ? 7'h1e : _T_183; // @[Mux.scala 47:69]
  wire [6:0] _T_185 = io_in[78] ? 7'h1d : _T_184; // @[Mux.scala 47:69]
  wire [6:0] _T_186 = io_in[79] ? 7'h1c : _T_185; // @[Mux.scala 47:69]
  wire [6:0] _T_187 = io_in[80] ? 7'h1b : _T_186; // @[Mux.scala 47:69]
  wire [6:0] _T_188 = io_in[81] ? 7'h1a : _T_187; // @[Mux.scala 47:69]
  wire [6:0] _T_189 = io_in[82] ? 7'h19 : _T_188; // @[Mux.scala 47:69]
  wire [6:0] _T_190 = io_in[83] ? 7'h18 : _T_189; // @[Mux.scala 47:69]
  wire [6:0] _T_191 = io_in[84] ? 7'h17 : _T_190; // @[Mux.scala 47:69]
  wire [6:0] _T_192 = io_in[85] ? 7'h16 : _T_191; // @[Mux.scala 47:69]
  wire [6:0] _T_193 = io_in[86] ? 7'h15 : _T_192; // @[Mux.scala 47:69]
  wire [6:0] _T_194 = io_in[87] ? 7'h14 : _T_193; // @[Mux.scala 47:69]
  wire [6:0] _T_195 = io_in[88] ? 7'h13 : _T_194; // @[Mux.scala 47:69]
  wire [6:0] _T_196 = io_in[89] ? 7'h12 : _T_195; // @[Mux.scala 47:69]
  wire [6:0] _T_197 = io_in[90] ? 7'h11 : _T_196; // @[Mux.scala 47:69]
  wire [6:0] _T_198 = io_in[91] ? 7'h10 : _T_197; // @[Mux.scala 47:69]
  wire [6:0] _T_199 = io_in[92] ? 7'hf : _T_198; // @[Mux.scala 47:69]
  wire [6:0] _T_200 = io_in[93] ? 7'he : _T_199; // @[Mux.scala 47:69]
  wire [6:0] _T_201 = io_in[94] ? 7'hd : _T_200; // @[Mux.scala 47:69]
  wire [6:0] _T_202 = io_in[95] ? 7'hc : _T_201; // @[Mux.scala 47:69]
  wire [6:0] _T_203 = io_in[96] ? 7'hb : _T_202; // @[Mux.scala 47:69]
  wire [6:0] _T_204 = io_in[97] ? 7'ha : _T_203; // @[Mux.scala 47:69]
  wire [6:0] _T_205 = io_in[98] ? 7'h9 : _T_204; // @[Mux.scala 47:69]
  wire [6:0] _T_206 = io_in[99] ? 7'h8 : _T_205; // @[Mux.scala 47:69]
  wire [6:0] _T_207 = io_in[100] ? 7'h7 : _T_206; // @[Mux.scala 47:69]
  wire [6:0] _T_208 = io_in[101] ? 7'h6 : _T_207; // @[Mux.scala 47:69]
  wire [6:0] _T_209 = io_in[102] ? 7'h5 : _T_208; // @[Mux.scala 47:69]
  wire [6:0] _T_210 = io_in[103] ? 7'h4 : _T_209; // @[Mux.scala 47:69]
  wire [6:0] _T_211 = io_in[104] ? 7'h3 : _T_210; // @[Mux.scala 47:69]
  wire [6:0] _T_212 = io_in[105] ? 7'h2 : _T_211; // @[Mux.scala 47:69]
  wire [6:0] _T_213 = io_in[106] ? 7'h1 : _T_212; // @[Mux.scala 47:69]
  assign io_out = io_in[107] ? 7'h0 : _T_213; // @[CLZ.scala 16:10]
endmodule
module RoundingUnit(
  input  [51:0] io_in,
  input         io_roundIn,
  input         io_stickyIn,
  input         io_signIn,
  input  [2:0]  io_rm,
  output [51:0] io_out,
  output        io_inexact,
  output        io_cout
);
  wire  g = io_in[0]; // @[RoundingUnit.scala 19:25]
  wire  inexact = io_roundIn | io_stickyIn; // @[RoundingUnit.scala 20:19]
  wire  _T_1 = io_roundIn & io_stickyIn; // @[RoundingUnit.scala 25:18]
  wire  _T_2 = ~io_stickyIn; // @[RoundingUnit.scala 25:33]
  wire  _T_3 = io_roundIn & _T_2; // @[RoundingUnit.scala 25:30]
  wire  _T_4 = _T_3 & g; // @[RoundingUnit.scala 25:36]
  wire  _T_5 = _T_1 | _T_4; // @[RoundingUnit.scala 25:24]
  wire  _T_6 = ~io_signIn; // @[RoundingUnit.scala 27:25]
  wire  _T_7 = inexact & _T_6; // @[RoundingUnit.scala 27:23]
  wire  _T_8 = inexact & io_signIn; // @[RoundingUnit.scala 28:23]
  wire  _T_9 = 3'h0 == io_rm; // @[Mux.scala 80:60]
  wire  _T_10 = _T_9 & _T_5; // @[Mux.scala 80:57]
  wire  _T_11 = 3'h1 == io_rm; // @[Mux.scala 80:60]
  wire  _T_12 = _T_11 ? 1'h0 : _T_10; // @[Mux.scala 80:57]
  wire  _T_13 = 3'h3 == io_rm; // @[Mux.scala 80:60]
  wire  _T_14 = _T_13 ? _T_7 : _T_12; // @[Mux.scala 80:57]
  wire  _T_15 = 3'h2 == io_rm; // @[Mux.scala 80:60]
  wire  _T_16 = _T_15 ? _T_8 : _T_14; // @[Mux.scala 80:57]
  wire  _T_17 = 3'h4 == io_rm; // @[Mux.scala 80:60]
  wire  r_up = _T_17 ? io_roundIn : _T_16; // @[Mux.scala 80:57]
  wire [51:0] out_r_up = io_in + 52'h1; // @[RoundingUnit.scala 32:24]
  wire  _T_20 = &io_in; // @[RoundingUnit.scala 36:28]
  assign io_out = r_up ? out_r_up : io_in; // @[RoundingUnit.scala 33:10]
  assign io_inexact = io_roundIn | io_stickyIn; // @[RoundingUnit.scala 34:14]
  assign io_cout = r_up & _T_20; // @[RoundingUnit.scala 36:11]
endmodule
module FMUL(
  input          clock,
  input          reset,
  input  [63:0]  io_a,
  input  [63:0]  io_b,
  input  [2:0]   io_rm,
  output [63:0]  io_result,
  output [4:0]   io_fflags,
  output         io_to_fadd_fp_prod_sign,
  output [10:0]  io_to_fadd_fp_prod_exp,
  output [104:0] io_to_fadd_fp_prod_sig,
  output         io_to_fadd_inter_flags_isNaN,
  output         io_to_fadd_inter_flags_isInf,
  output         io_to_fadd_inter_flags_isInv,
  output         io_to_fadd_inter_flags_overflow
);
  wire [107:0] CLZ_io_in; // @[CLZ.scala 21:21]
  wire [6:0] CLZ_io_out; // @[CLZ.scala 21:21]
  wire [51:0] tininess_rounder_io_in; // @[RoundingUnit.scala 44:25]
  wire  tininess_rounder_io_roundIn; // @[RoundingUnit.scala 44:25]
  wire  tininess_rounder_io_stickyIn; // @[RoundingUnit.scala 44:25]
  wire  tininess_rounder_io_signIn; // @[RoundingUnit.scala 44:25]
  wire [2:0] tininess_rounder_io_rm; // @[RoundingUnit.scala 44:25]
  wire [51:0] tininess_rounder_io_out; // @[RoundingUnit.scala 44:25]
  wire  tininess_rounder_io_inexact; // @[RoundingUnit.scala 44:25]
  wire  tininess_rounder_io_cout; // @[RoundingUnit.scala 44:25]
  wire [51:0] rounder_io_in; // @[RoundingUnit.scala 44:25]
  wire  rounder_io_roundIn; // @[RoundingUnit.scala 44:25]
  wire  rounder_io_stickyIn; // @[RoundingUnit.scala 44:25]
  wire  rounder_io_signIn; // @[RoundingUnit.scala 44:25]
  wire [2:0] rounder_io_rm; // @[RoundingUnit.scala 44:25]
  wire [51:0] rounder_io_out; // @[RoundingUnit.scala 44:25]
  wire  rounder_io_inexact; // @[RoundingUnit.scala 44:25]
  wire  rounder_io_cout; // @[RoundingUnit.scala 44:25]
  wire  fp_a_sign = io_a[63]; // @[package.scala 59:19]
  wire [10:0] fp_a_exp = io_a[62:52]; // @[package.scala 60:18]
  wire [51:0] fp_a_sig = io_a[51:0]; // @[package.scala 61:18]
  wire  fp_b_sign = io_b[63]; // @[package.scala 59:19]
  wire [10:0] fp_b_exp = io_b[62:52]; // @[package.scala 60:18]
  wire [51:0] fp_b_sig = io_b[51:0]; // @[package.scala 61:18]
  wire  decode_a_expNotZero = |fp_a_exp; // @[package.scala 32:28]
  wire  decode_a_expIsOnes = &fp_a_exp; // @[package.scala 33:27]
  wire  decode_a_sigNotZero = |fp_a_sig; // @[package.scala 34:28]
  wire  decode_a_expIsZero = ~decode_a_expNotZero; // @[package.scala 37:27]
  wire  decode_a_sigIsZero = ~decode_a_sigNotZero; // @[package.scala 40:27]
  wire  decode_a_isInf = decode_a_expIsOnes & decode_a_sigIsZero; // @[package.scala 42:40]
  wire  decode_a_isZero = decode_a_expIsZero & decode_a_sigIsZero; // @[package.scala 43:41]
  wire  decode_a_isNaN = decode_a_expIsOnes & decode_a_sigNotZero; // @[package.scala 44:40]
  wire  _T_17 = ~fp_a_sig[51]; // @[package.scala 45:40]
  wire  decode_a_isSNaN = decode_a_isNaN & _T_17; // @[package.scala 45:37]
  wire  decode_b_expNotZero = |fp_b_exp; // @[package.scala 32:28]
  wire  decode_b_expIsOnes = &fp_b_exp; // @[package.scala 33:27]
  wire  decode_b_sigNotZero = |fp_b_sig; // @[package.scala 34:28]
  wire  decode_b_expIsZero = ~decode_b_expNotZero; // @[package.scala 37:27]
  wire  decode_b_sigIsZero = ~decode_b_sigNotZero; // @[package.scala 40:27]
  wire  decode_b_isInf = decode_b_expIsOnes & decode_b_sigIsZero; // @[package.scala 42:40]
  wire  decode_b_isZero = decode_b_expIsZero & decode_b_sigIsZero; // @[package.scala 43:41]
  wire  decode_b_isNaN = decode_b_expIsOnes & decode_b_sigNotZero; // @[package.scala 44:40]
  wire  _T_33 = ~fp_b_sig[51]; // @[package.scala 45:40]
  wire  decode_b_isSNaN = decode_b_isNaN & _T_33; // @[package.scala 45:37]
  wire [10:0] _GEN_0 = {{10'd0}, decode_a_expIsZero}; // @[package.scala 83:27]
  wire [10:0] raw_a_exp = fp_a_exp | _GEN_0; // @[package.scala 83:27]
  wire [52:0] raw_a_sig = {decode_a_expNotZero,fp_a_sig}; // @[Cat.scala 29:58]
  wire [10:0] _GEN_1 = {{10'd0}, decode_b_expIsZero}; // @[package.scala 83:27]
  wire [10:0] raw_b_exp = fp_b_exp | _GEN_1; // @[package.scala 83:27]
  wire [52:0] raw_b_sig = {decode_b_expNotZero,fp_b_sig}; // @[Cat.scala 29:58]
  wire  prod_sign = fp_a_sign ^ fp_b_sign; // @[FMUL.scala 35:29]
  wire [11:0] exp_sum = raw_a_exp + raw_b_exp; // @[FMUL.scala 52:27]
  wire [11:0] prod_exp = exp_sum - 12'h3c7; // @[FMUL.scala 53:26]
  wire [12:0] _T_45 = {1'h0,exp_sum}; // @[Cat.scala 29:58]
  wire [12:0] shift_lim_sub = _T_45 - 13'h3c8; // @[FMUL.scala 55:46]
  wire  prod_exp_uf = shift_lim_sub[12]; // @[FMUL.scala 56:39]
  wire [11:0] shift_lim = shift_lim_sub[11:0]; // @[FMUL.scala 57:37]
  wire  prod_exp_ov = exp_sum > 12'hbfd; // @[FMUL.scala 59:29]
  wire [52:0] subnormal_sig = decode_a_expIsZero ? raw_a_sig : raw_b_sig; // @[FMUL.scala 62:26]
  wire [11:0] _GEN_2 = {{5'd0}, CLZ_io_out}; // @[FMUL.scala 64:30]
  wire  exceed_lim = shift_lim <= _GEN_2; // @[FMUL.scala 64:30]
  wire [11:0] _T_49 = exceed_lim ? shift_lim : {{5'd0}, CLZ_io_out}; // @[FMUL.scala 65:44]
  wire [11:0] shift_amt = prod_exp_uf ? 12'h0 : _T_49; // @[FMUL.scala 65:22]
  wire [105:0] prod = raw_a_sig * raw_b_sig; // @[FMUL.scala 67:24]
  wire [160:0] sig_shifter_in = {55'h0,prod}; // @[Cat.scala 29:58]
  wire [4255:0] _GEN_3 = {{4095'd0}, sig_shifter_in}; // @[FMUL.scala 69:41]
  wire [4255:0] _T_50 = _GEN_3 << shift_amt; // @[FMUL.scala 69:41]
  wire [160:0] sig_shifted_raw = _T_50[160:0]; // @[FMUL.scala 69:54]
  wire [11:0] exp_shifted = prod_exp - shift_amt; // @[FMUL.scala 70:30]
  wire  _T_52 = exceed_lim | prod_exp_uf; // @[FMUL.scala 71:38]
  wire  _T_55 = ~sig_shifted_raw[160]; // @[FMUL.scala 71:57]
  wire  exp_is_subnormal = _T_52 & _T_55; // @[FMUL.scala 71:54]
  wire  no_extra_shift = sig_shifted_raw[160] | exp_is_subnormal; // @[FMUL.scala 72:55]
  wire [11:0] _T_59 = exp_shifted - 12'h1; // @[FMUL.scala 74:95]
  wire [11:0] _T_60 = no_extra_shift ? exp_shifted : _T_59; // @[FMUL.scala 74:53]
  wire [11:0] exp_pre_round = exp_is_subnormal ? 12'h0 : _T_60; // @[FMUL.scala 74:26]
  wire [160:0] _T_62 = {sig_shifted_raw[159:0],1'h0}; // @[Cat.scala 29:58]
  wire [160:0] sig_shifted = no_extra_shift ? sig_shifted_raw : _T_62; // @[FMUL.scala 75:24]
  wire  _T_71 = sig_shifted[160:159] == 2'h0; // @[FMUL.scala 84:38]
  wire  _T_73 = sig_shifted[160:159] == 2'h1; // @[FMUL.scala 85:26]
  wire  _T_74 = ~tininess_rounder_io_cout; // @[FMUL.scala 85:46]
  wire  _T_75 = _T_73 & _T_74; // @[FMUL.scala 85:43]
  wire  tininess = _T_71 | _T_75; // @[FMUL.scala 84:55]
  wire [11:0] _GEN_4 = {{11'd0}, rounder_io_cout}; // @[FMUL.scala 94:37]
  wire [11:0] exp_rounded = _GEN_4 + exp_pre_round; // @[FMUL.scala 94:37]
  wire  _T_84 = exp_pre_round == 12'h7fe; // @[FMUL.scala 99:19]
  wire  _T_85 = exp_pre_round == 12'h7ff; // @[FMUL.scala 100:19]
  wire  _T_86 = rounder_io_cout ? _T_84 : _T_85; // @[FMUL.scala 97:22]
  wire  common_of = _T_86 | prod_exp_ov; // @[FMUL.scala 101:5]
  wire  common_ix = rounder_io_inexact | common_of; // @[FMUL.scala 102:38]
  wire  common_uf = tininess & common_ix; // @[FMUL.scala 103:28]
  wire  _T_87 = io_rm == 3'h1; // @[RoundingUnit.scala 54:8]
  wire  _T_88 = io_rm == 3'h2; // @[RoundingUnit.scala 54:23]
  wire  _T_89 = ~prod_sign; // @[RoundingUnit.scala 54:34]
  wire  _T_90 = _T_88 & _T_89; // @[RoundingUnit.scala 54:31]
  wire  _T_91 = _T_87 | _T_90; // @[RoundingUnit.scala 54:16]
  wire  _T_92 = io_rm == 3'h3; // @[RoundingUnit.scala 54:48]
  wire  _T_93 = _T_92 & prod_sign; // @[RoundingUnit.scala 54:56]
  wire  rmin = _T_91 | _T_93; // @[RoundingUnit.scala 54:41]
  wire [10:0] of_exp = rmin ? 11'h7fe : 11'h7ff; // @[FMUL.scala 107:19]
  wire [10:0] common_exp = common_of ? of_exp : exp_rounded[10:0]; // @[FMUL.scala 111:23]
  wire [51:0] _T_96 = rmin ? 52'hfffffffffffff : 52'h0; // @[FMUL.scala 118:8]
  wire [51:0] common_sig = common_of ? _T_96 : rounder_io_out; // @[FMUL.scala 116:23]
  wire [63:0] common_result = {prod_sign,common_exp,common_sig}; // @[Cat.scala 29:58]
  wire [4:0] common_fflags = {2'h0,common_of,common_uf,common_ix}; // @[Cat.scala 29:58]
  wire  hasZero = decode_a_isZero | decode_b_isZero; // @[FMUL.scala 129:33]
  wire  hasNaN = decode_a_isNaN | decode_b_isNaN; // @[FMUL.scala 130:31]
  wire  hasSNaN = decode_a_isSNaN | decode_b_isSNaN; // @[FMUL.scala 131:33]
  wire  hasInf = decode_a_isInf | decode_b_isInf; // @[FMUL.scala 132:31]
  wire  _T_101 = hasZero | hasNaN; // @[FMUL.scala 133:37]
  wire  special_case_happen = _T_101 | hasInf; // @[FMUL.scala 133:47]
  wire  zero_mul_inf = hasZero & hasInf; // @[FMUL.scala 135:30]
  wire  nan_result = hasNaN | zero_mul_inf; // @[FMUL.scala 136:27]
  wire  special_iv = hasSNaN | zero_mul_inf; // @[FMUL.scala 140:28]
  wire [63:0] _T_108 = {prod_sign,11'h7ff,52'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_109 = {prod_sign,63'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_110 = hasInf ? _T_108 : _T_109; // @[FMUL.scala 145:8]
  wire [63:0] special_result = nan_result ? 64'h7ff8000000000000 : _T_110; // @[FMUL.scala 143:27]
  wire [4:0] special_fflags = {special_iv,1'h0,1'h0,2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_116 = hasZero ? 12'h0 : exp_pre_round; // @[FMUL.scala 156:32]
  wire  _T_120 = |sig_shifted[54:0]; // @[FMUL.scala 159:83]
  wire [104:0] _GEN_5 = {{104'd0}, _T_120}; // @[FMUL.scala 159:49]
  wire [104:0] _T_121 = sig_shifted[159:55] | _GEN_5; // @[FMUL.scala 159:49]
  wire  _T_123 = ~nan_result; // @[FMUL.scala 162:45]
  CLZ CLZ ( // @[CLZ.scala 21:21]
    .io_in(CLZ_io_in),
    .io_out(CLZ_io_out)
  );
  RoundingUnit tininess_rounder ( // @[RoundingUnit.scala 44:25]
    .io_in(tininess_rounder_io_in),
    .io_roundIn(tininess_rounder_io_roundIn),
    .io_stickyIn(tininess_rounder_io_stickyIn),
    .io_signIn(tininess_rounder_io_signIn),
    .io_rm(tininess_rounder_io_rm),
    .io_out(tininess_rounder_io_out),
    .io_inexact(tininess_rounder_io_inexact),
    .io_cout(tininess_rounder_io_cout)
  );
  RoundingUnit rounder ( // @[RoundingUnit.scala 44:25]
    .io_in(rounder_io_in),
    .io_roundIn(rounder_io_roundIn),
    .io_stickyIn(rounder_io_stickyIn),
    .io_signIn(rounder_io_signIn),
    .io_rm(rounder_io_rm),
    .io_out(rounder_io_out),
    .io_inexact(rounder_io_inexact),
    .io_cout(rounder_io_cout)
  );
  assign io_result = special_case_happen ? special_result : common_result; // @[FMUL.scala 152:13]
  assign io_fflags = special_case_happen ? special_fflags : common_fflags; // @[FMUL.scala 153:13]
  assign io_to_fadd_fp_prod_sign = fp_a_sign ^ fp_b_sign; // @[FMUL.scala 155:27]
  assign io_to_fadd_fp_prod_exp = _T_116[10:0]; // @[FMUL.scala 156:26]
  assign io_to_fadd_fp_prod_sig = hasZero ? 105'h0 : _T_121; // @[FMUL.scala 157:26]
  assign io_to_fadd_inter_flags_isNaN = hasNaN | zero_mul_inf; // @[FMUL.scala 163:32]
  assign io_to_fadd_inter_flags_isInf = hasInf & _T_123; // @[FMUL.scala 162:32]
  assign io_to_fadd_inter_flags_isInv = hasSNaN | zero_mul_inf; // @[FMUL.scala 161:32]
  assign io_to_fadd_inter_flags_overflow = exp_pre_round > 12'h7ff; // @[FMUL.scala 164:35]
  assign CLZ_io_in = {55'h0,subnormal_sig}; // @[CLZ.scala 22:15]
  assign tininess_rounder_io_in = sig_shifted[158:107]; // @[RoundingUnit.scala 45:19]
  assign tininess_rounder_io_roundIn = sig_shifted[106]; // @[RoundingUnit.scala 46:24]
  assign tininess_rounder_io_stickyIn = |sig_shifted[105:0]; // @[RoundingUnit.scala 47:25]
  assign tininess_rounder_io_signIn = fp_a_sign ^ fp_b_sign; // @[RoundingUnit.scala 49:23]
  assign tininess_rounder_io_rm = io_rm; // @[RoundingUnit.scala 48:19]
  assign rounder_io_in = sig_shifted[159:108]; // @[RoundingUnit.scala 45:19]
  assign rounder_io_roundIn = sig_shifted[107]; // @[RoundingUnit.scala 46:24]
  assign rounder_io_stickyIn = |sig_shifted[106:0]; // @[RoundingUnit.scala 47:25]
  assign rounder_io_signIn = fp_a_sign ^ fp_b_sign; // @[RoundingUnit.scala 49:23]
  assign rounder_io_rm = io_rm; // @[RoundingUnit.scala 48:19]
endmodule
