module MultiDimTime(
  input         clock,
  input         reset,
  input         io_in,
  output [1:0]  io_out_0,
  output [1:0]  io_out_1,
  output [1:0]  io_out_2,
  output [1:0]  io_out_3,
  output [1:0]  io_out_4,
  output [17:0] io_index_0,
  output [17:0] io_index_1,
  output [17:0] io_index_2,
  output [17:0] io_index_3
);
  reg [15:0] regs_0; // @[mem.scala 81:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 81:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 81:12]
  reg [31:0] _RAND_2;
  reg [15:0] regs_3; // @[mem.scala 81:12]
  reg [31:0] _RAND_3;
  reg [15:0] regs_4; // @[mem.scala 81:12]
  reg [31:0] _RAND_4;
  wire [15:0] _GEN_10 = {{15'd0}, io_in}; // @[mem.scala 95:42]
  wire [15:0] _T_1 = regs_0 + _GEN_10; // @[mem.scala 95:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 95:48]
  wire [15:0] _T_3 = regs_1 + _GEN_10; // @[mem.scala 95:42]
  wire  back_1 = _T_3 == 16'h14; // @[mem.scala 95:48]
  wire [15:0] _T_5 = regs_2 + _GEN_10; // @[mem.scala 95:42]
  wire  back_2 = _T_5 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_7 = regs_3 + _GEN_10; // @[mem.scala 95:42]
  wire  back_3 = _T_7 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_9 = regs_4 + _GEN_10; // @[mem.scala 95:42]
  wire  back_4 = _T_9 == 16'h6; // @[mem.scala 95:48]
  wire  _T_10 = ~back_0; // @[mem.scala 102:20]
  wire [1:0] _T_11 = {_T_10, 1'h0}; // @[mem.scala 102:31]
  wire  _T_12 = ~back_1; // @[mem.scala 102:40]
  wire [1:0] _GEN_15 = {{1'd0}, _T_12}; // @[mem.scala 102:37]
  wire  _T_16 = back_0 & back_1; // @[mem.scala 101:46]
  wire  _T_17 = ~_T_16; // @[mem.scala 102:20]
  wire [1:0] _T_18 = {_T_17, 1'h0}; // @[mem.scala 102:31]
  wire  _T_19 = ~back_2; // @[mem.scala 102:40]
  wire [1:0] _GEN_17 = {{1'd0}, _T_19}; // @[mem.scala 102:37]
  wire  _T_24 = _T_16 & back_2; // @[mem.scala 101:46]
  wire  _T_25 = ~_T_24; // @[mem.scala 102:20]
  wire [1:0] _T_26 = {_T_25, 1'h0}; // @[mem.scala 102:31]
  wire  _T_27 = ~back_3; // @[mem.scala 102:40]
  wire [1:0] _GEN_19 = {{1'd0}, _T_27}; // @[mem.scala 102:37]
  wire  _T_33 = _T_24 & back_3; // @[mem.scala 101:46]
  wire  _T_34 = ~_T_33; // @[mem.scala 102:20]
  wire [1:0] _T_35 = {_T_34, 1'h0}; // @[mem.scala 102:31]
  wire  _T_36 = ~back_4; // @[mem.scala 102:40]
  wire [1:0] _GEN_21 = {{1'd0}, _T_36}; // @[mem.scala 102:37]
  wire  _GEN_9 = back_0 ? 1'h0 : io_in; // @[mem.scala 112:16]
  assign io_out_0 = {{1'd0}, _GEN_9}; // @[mem.scala 114:15 mem.scala 117:15]
  assign io_out_1 = _T_11 | _GEN_15; // @[mem.scala 102:15]
  assign io_out_2 = _T_18 | _GEN_17; // @[mem.scala 102:15]
  assign io_out_3 = _T_26 | _GEN_19; // @[mem.scala 102:15]
  assign io_out_4 = _T_35 | _GEN_21; // @[mem.scala 102:15]
  assign io_index_0 = {{2'd0}, regs_0}; // @[mem.scala 111:15]
  assign io_index_1 = {{2'd0}, regs_1}; // @[mem.scala 99:17]
  assign io_index_2 = {{2'd0}, regs_2}; // @[mem.scala 99:17]
  assign io_index_3 = {{2'd0}, regs_3}; // @[mem.scala 99:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (_T_16) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
    if (reset) begin
      regs_3 <= 16'h0;
    end else if (_T_24) begin
      if (back_3) begin
        regs_3 <= 16'h0;
      end else begin
        regs_3 <= _T_7;
      end
    end
    if (reset) begin
      regs_4 <= 16'h0;
    end else if (_T_33) begin
      if (back_4) begin
        regs_4 <= 16'h0;
      end else begin
        regs_4 <= _T_9;
      end
    end
  end
endmodule
module ComputeCell_Latency(
  input         clock,
  input         reset,
  input  [15:0] io_data_2_in,
  input  [15:0] io_data_1_in,
  input  [15:0] io_data_0_in,
  output [15:0] io_data_0_out
);
  reg [15:0] _T_4_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_0;
  reg [15:0] _T_5_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  reg [15:0] _T_6_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [15:0] _T_7_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [15:0] _T_8_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [15:0] _T_9_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [15:0] _T_10_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [15:0] _T_11_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [15:0] _T_12_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  reg [15:0] _T_13_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_9;
  reg [15:0] _T_14_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_10;
  reg [15:0] delay_a_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg [15:0] _T_16_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg [15:0] _T_17_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg [15:0] _T_18_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  reg [15:0] _T_19_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  reg [15:0] _T_20_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg [15:0] _T_21_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  reg [15:0] _T_22_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_18;
  reg [15:0] _T_23_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_19;
  reg [15:0] _T_24_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_20;
  reg [15:0] _T_25_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_21;
  reg [15:0] _T_26_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_22;
  reg [15:0] delay_b_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_23;
  reg [15:0] _T_28_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_24;
  reg [15:0] _T_29_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_25;
  reg [15:0] _T_30_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_26;
  reg [15:0] _T_31_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_27;
  reg [15:0] _T_32_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_28;
  reg [15:0] _T_33_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_29;
  reg [15:0] _T_34_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_30;
  reg [15:0] _T_35_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_31;
  reg [15:0] _T_36_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_32;
  reg [15:0] _T_37_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_33;
  reg [15:0] _T_38_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_34;
  reg [15:0] delay_c_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_35;
  wire [31:0] _T_42 = delay_a_0 * delay_b_0; // @[cell.scala 145:63]
  wire [31:0] _GEN_36 = {{16'd0}, delay_c_0}; // @[cell.scala 145:50]
  wire [31:0] _T_44 = _GEN_36 + _T_42; // @[cell.scala 145:50]
  assign io_data_0_out = _T_44[15:0]; // @[cell.scala 148:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_5_0 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_6_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_7_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_8_0 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_9_0 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_10_0 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_11_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_12_0 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_13_0 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_14_0 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  delay_a_0 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_16_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_17_0 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_18_0 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_19_0 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_20_0 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_21_0 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_22_0 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_23_0 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_24_0 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_25_0 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_26_0 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  delay_b_0 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_28_0 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_29_0 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_30_0 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_31_0 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_32_0 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_33_0 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_34_0 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_35_0 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_36_0 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_37_0 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_38_0 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  delay_c_0 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_4_0 <= 16'h0;
    end else begin
      _T_4_0 <= io_data_1_in;
    end
    if (reset) begin
      _T_5_0 <= 16'h0;
    end else begin
      _T_5_0 <= _T_4_0;
    end
    if (reset) begin
      _T_6_0 <= 16'h0;
    end else begin
      _T_6_0 <= _T_5_0;
    end
    if (reset) begin
      _T_7_0 <= 16'h0;
    end else begin
      _T_7_0 <= _T_6_0;
    end
    if (reset) begin
      _T_8_0 <= 16'h0;
    end else begin
      _T_8_0 <= _T_7_0;
    end
    if (reset) begin
      _T_9_0 <= 16'h0;
    end else begin
      _T_9_0 <= _T_8_0;
    end
    if (reset) begin
      _T_10_0 <= 16'h0;
    end else begin
      _T_10_0 <= _T_9_0;
    end
    if (reset) begin
      _T_11_0 <= 16'h0;
    end else begin
      _T_11_0 <= _T_10_0;
    end
    if (reset) begin
      _T_12_0 <= 16'h0;
    end else begin
      _T_12_0 <= _T_11_0;
    end
    if (reset) begin
      _T_13_0 <= 16'h0;
    end else begin
      _T_13_0 <= _T_12_0;
    end
    if (reset) begin
      _T_14_0 <= 16'h0;
    end else begin
      _T_14_0 <= _T_13_0;
    end
    if (reset) begin
      delay_a_0 <= 16'h0;
    end else begin
      delay_a_0 <= _T_14_0;
    end
    if (reset) begin
      _T_16_0 <= 16'h0;
    end else begin
      _T_16_0 <= io_data_2_in;
    end
    if (reset) begin
      _T_17_0 <= 16'h0;
    end else begin
      _T_17_0 <= _T_16_0;
    end
    if (reset) begin
      _T_18_0 <= 16'h0;
    end else begin
      _T_18_0 <= _T_17_0;
    end
    if (reset) begin
      _T_19_0 <= 16'h0;
    end else begin
      _T_19_0 <= _T_18_0;
    end
    if (reset) begin
      _T_20_0 <= 16'h0;
    end else begin
      _T_20_0 <= _T_19_0;
    end
    if (reset) begin
      _T_21_0 <= 16'h0;
    end else begin
      _T_21_0 <= _T_20_0;
    end
    if (reset) begin
      _T_22_0 <= 16'h0;
    end else begin
      _T_22_0 <= _T_21_0;
    end
    if (reset) begin
      _T_23_0 <= 16'h0;
    end else begin
      _T_23_0 <= _T_22_0;
    end
    if (reset) begin
      _T_24_0 <= 16'h0;
    end else begin
      _T_24_0 <= _T_23_0;
    end
    if (reset) begin
      _T_25_0 <= 16'h0;
    end else begin
      _T_25_0 <= _T_24_0;
    end
    if (reset) begin
      _T_26_0 <= 16'h0;
    end else begin
      _T_26_0 <= _T_25_0;
    end
    if (reset) begin
      delay_b_0 <= 16'h0;
    end else begin
      delay_b_0 <= _T_26_0;
    end
    if (reset) begin
      _T_28_0 <= 16'h0;
    end else begin
      _T_28_0 <= io_data_0_in;
    end
    if (reset) begin
      _T_29_0 <= 16'h0;
    end else begin
      _T_29_0 <= _T_28_0;
    end
    if (reset) begin
      _T_30_0 <= 16'h0;
    end else begin
      _T_30_0 <= _T_29_0;
    end
    if (reset) begin
      _T_31_0 <= 16'h0;
    end else begin
      _T_31_0 <= _T_30_0;
    end
    if (reset) begin
      _T_32_0 <= 16'h0;
    end else begin
      _T_32_0 <= _T_31_0;
    end
    if (reset) begin
      _T_33_0 <= 16'h0;
    end else begin
      _T_33_0 <= _T_32_0;
    end
    if (reset) begin
      _T_34_0 <= 16'h0;
    end else begin
      _T_34_0 <= _T_33_0;
    end
    if (reset) begin
      _T_35_0 <= 16'h0;
    end else begin
      _T_35_0 <= _T_34_0;
    end
    if (reset) begin
      _T_36_0 <= 16'h0;
    end else begin
      _T_36_0 <= _T_35_0;
    end
    if (reset) begin
      _T_37_0 <= 16'h0;
    end else begin
      _T_37_0 <= _T_36_0;
    end
    if (reset) begin
      _T_38_0 <= 16'h0;
    end else begin
      _T_38_0 <= _T_37_0;
    end
    if (reset) begin
      delay_c_0 <= 16'h0;
    end else begin
      delay_c_0 <= _T_38_0;
    end
  end
endmodule
module SystolicOutput(
  input         io_port_in_valid,
  input  [15:0] io_port_in_bits,
  output        io_port_out_valid,
  output [15:0] io_port_out_bits,
  input         io_from_cell_valid,
  input  [15:0] io_from_cell_bits,
  output        io_to_cell_valid,
  output [15:0] io_to_cell_bits
);
  assign io_port_out_valid = io_from_cell_valid; // @[pe_modules.scala 111:15]
  assign io_port_out_bits = io_from_cell_bits; // @[pe_modules.scala 111:15]
  assign io_to_cell_valid = io_port_in_valid; // @[pe_modules.scala 110:14]
  assign io_to_cell_bits = io_port_in_bits; // @[pe_modules.scala 110:14]
endmodule
module StationaryInput_Pipeline(
  input         clock,
  input         reset,
  input         io_port_in_valid,
  input  [15:0] io_port_in_bits,
  output        io_port_out_valid,
  output [15:0] io_port_out_bits,
  output [15:0] io_to_cell_bits,
  input         io_sig_stat2trans
);
  reg  trans_valid; // @[pe_modules.scala 128:22]
  reg [31:0] _RAND_0;
  reg [15:0] trans_bits; // @[pe_modules.scala 128:22]
  reg [31:0] _RAND_1;
  reg  update_valid; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_2;
  reg [15:0] update_bits_0; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_3;
  reg [15:0] update_bits_1; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_4;
  reg [15:0] update_bits_2; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_5;
  reg [15:0] update_bits_3; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_6;
  reg [15:0] update_bits_4; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_7;
  reg [15:0] update_bits_5; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_8;
  reg [15:0] update_bits_6; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_9;
  reg [15:0] update_bits_7; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_10;
  reg [15:0] update_bits_8; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_11;
  reg [15:0] update_bits_9; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_12;
  reg [15:0] update_bits_10; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_13;
  reg [15:0] update_bits_11; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_14;
  reg  stat_valid; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_15;
  reg [15:0] stat_bits_0; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_16;
  reg [15:0] stat_bits_1; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_17;
  reg [15:0] stat_bits_2; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_18;
  reg [15:0] stat_bits_3; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_19;
  reg [15:0] stat_bits_4; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_20;
  reg [15:0] stat_bits_5; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_21;
  reg [15:0] stat_bits_6; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_22;
  reg [15:0] stat_bits_7; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_23;
  reg [15:0] stat_bits_8; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_24;
  reg [15:0] stat_bits_9; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_25;
  reg [15:0] stat_bits_10; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_26;
  reg [15:0] stat_bits_11; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_27;
  reg  reg_stat2trans_0; // @[pe_modules.scala 135:31]
  reg [31:0] _RAND_28;
  reg [3:0] write_trans_pos; // @[pe_modules.scala 137:32]
  reg [31:0] _RAND_29;
  reg [3:0] read_stat_pos; // @[pe_modules.scala 138:30]
  reg [31:0] _RAND_30;
  wire  _T_4 = ~update_valid; // @[pe_modules.scala 142:26]
  wire [3:0] _GEN_51 = {{3'd0}, trans_valid}; // @[pe_modules.scala 142:60]
  wire [3:0] _T_6 = write_trans_pos + _GEN_51; // @[pe_modules.scala 142:60]
  wire  _T_7 = _T_6 == 4'hc; // @[pe_modules.scala 142:79]
  wire  _T_13 = _T_4 & trans_valid; // @[pe_modules.scala 143:24]
  wire [3:0] _T_15 = read_stat_pos + 4'h1; // @[pe_modules.scala 148:53]
  wire  _T_16 = _T_15 == 4'hc; // @[pe_modules.scala 148:57]
  wire  _T_21 = write_trans_pos == 4'hb; // @[pe_modules.scala 149:23]
  wire  _T_22 = _T_21 & trans_valid; // @[pe_modules.scala 149:45]
  wire  _GEN_24 = _T_22 | update_valid; // @[pe_modules.scala 149:60]
  reg [15:0] _T_24; // @[pe_modules.scala 163:29]
  reg [31:0] _RAND_31;
  assign io_port_out_valid = update_valid; // @[pe_modules.scala 139:21]
  assign io_port_out_bits = trans_bits; // @[pe_modules.scala 140:20]
  assign io_to_cell_bits = _T_24; // @[pe_modules.scala 163:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  trans_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  trans_bits = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  update_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  update_bits_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  update_bits_1 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  update_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  update_bits_3 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  update_bits_4 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  update_bits_5 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  update_bits_6 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  update_bits_7 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  update_bits_8 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  update_bits_9 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  update_bits_10 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  update_bits_11 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  stat_valid = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  stat_bits_0 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  stat_bits_1 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  stat_bits_2 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  stat_bits_3 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  stat_bits_4 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  stat_bits_5 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  stat_bits_6 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  stat_bits_7 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  stat_bits_8 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  stat_bits_9 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  stat_bits_10 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  stat_bits_11 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  reg_stat2trans_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  write_trans_pos = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  read_stat_pos = _RAND_30[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_24 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      trans_valid <= 1'h0;
    end else begin
      trans_valid <= io_port_in_valid;
    end
    if (reset) begin
      trans_bits <= 16'h0;
    end else begin
      trans_bits <= io_port_in_bits;
    end
    if (reset) begin
      update_valid <= 1'h0;
    end else if (reg_stat2trans_0) begin
      update_valid <= 1'h0;
    end else begin
      update_valid <= _GEN_24;
    end
    if (reset) begin
      update_bits_0 <= 16'h0;
    end else if (_T_13) begin
      if (4'h0 == write_trans_pos) begin
        update_bits_0 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_1 <= 16'h0;
    end else if (_T_13) begin
      if (4'h1 == write_trans_pos) begin
        update_bits_1 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_2 <= 16'h0;
    end else if (_T_13) begin
      if (4'h2 == write_trans_pos) begin
        update_bits_2 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_3 <= 16'h0;
    end else if (_T_13) begin
      if (4'h3 == write_trans_pos) begin
        update_bits_3 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_4 <= 16'h0;
    end else if (_T_13) begin
      if (4'h4 == write_trans_pos) begin
        update_bits_4 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_5 <= 16'h0;
    end else if (_T_13) begin
      if (4'h5 == write_trans_pos) begin
        update_bits_5 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_6 <= 16'h0;
    end else if (_T_13) begin
      if (4'h6 == write_trans_pos) begin
        update_bits_6 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_7 <= 16'h0;
    end else if (_T_13) begin
      if (4'h7 == write_trans_pos) begin
        update_bits_7 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_8 <= 16'h0;
    end else if (_T_13) begin
      if (4'h8 == write_trans_pos) begin
        update_bits_8 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_9 <= 16'h0;
    end else if (_T_13) begin
      if (4'h9 == write_trans_pos) begin
        update_bits_9 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_10 <= 16'h0;
    end else if (_T_13) begin
      if (4'ha == write_trans_pos) begin
        update_bits_10 <= trans_bits;
      end
    end
    if (reset) begin
      update_bits_11 <= 16'h0;
    end else if (_T_13) begin
      if (4'hb == write_trans_pos) begin
        update_bits_11 <= trans_bits;
      end
    end
    if (reset) begin
      stat_valid <= 1'h0;
    end else if (reg_stat2trans_0) begin
      stat_valid <= update_valid;
    end
    if (reset) begin
      stat_bits_0 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_0 <= update_bits_0;
    end
    if (reset) begin
      stat_bits_1 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_1 <= update_bits_1;
    end
    if (reset) begin
      stat_bits_2 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_2 <= update_bits_2;
    end
    if (reset) begin
      stat_bits_3 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_3 <= update_bits_3;
    end
    if (reset) begin
      stat_bits_4 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_4 <= update_bits_4;
    end
    if (reset) begin
      stat_bits_5 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_5 <= update_bits_5;
    end
    if (reset) begin
      stat_bits_6 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_6 <= update_bits_6;
    end
    if (reset) begin
      stat_bits_7 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_7 <= update_bits_7;
    end
    if (reset) begin
      stat_bits_8 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_8 <= update_bits_8;
    end
    if (reset) begin
      stat_bits_9 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_9 <= update_bits_9;
    end
    if (reset) begin
      stat_bits_10 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_10 <= update_bits_10;
    end
    if (reset) begin
      stat_bits_11 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_11 <= update_bits_11;
    end
    if (reset) begin
      reg_stat2trans_0 <= 1'h0;
    end else begin
      reg_stat2trans_0 <= io_sig_stat2trans;
    end
    if (reset) begin
      write_trans_pos <= 4'h0;
    end else if (_T_4) begin
      if (_T_7) begin
        write_trans_pos <= 4'h0;
      end else begin
        write_trans_pos <= _T_6;
      end
    end
    if (reset) begin
      read_stat_pos <= 4'h0;
    end else if (stat_valid) begin
      if (_T_16) begin
        read_stat_pos <= 4'h0;
      end else begin
        read_stat_pos <= _T_15;
      end
    end
    if (reset) begin
      _T_24 <= 16'h0;
    end else if (4'hb == read_stat_pos) begin
      _T_24 <= stat_bits_11;
    end else if (4'ha == read_stat_pos) begin
      _T_24 <= stat_bits_10;
    end else if (4'h9 == read_stat_pos) begin
      _T_24 <= stat_bits_9;
    end else if (4'h8 == read_stat_pos) begin
      _T_24 <= stat_bits_8;
    end else if (4'h7 == read_stat_pos) begin
      _T_24 <= stat_bits_7;
    end else if (4'h6 == read_stat_pos) begin
      _T_24 <= stat_bits_6;
    end else if (4'h5 == read_stat_pos) begin
      _T_24 <= stat_bits_5;
    end else if (4'h4 == read_stat_pos) begin
      _T_24 <= stat_bits_4;
    end else if (4'h3 == read_stat_pos) begin
      _T_24 <= stat_bits_3;
    end else if (4'h2 == read_stat_pos) begin
      _T_24 <= stat_bits_2;
    end else if (4'h1 == read_stat_pos) begin
      _T_24 <= stat_bits_1;
    end else begin
      _T_24 <= stat_bits_0;
    end
  end
endmodule
module SystolicInput(
  input         clock,
  input         reset,
  input         io_port_in_valid,
  input  [15:0] io_port_in_bits,
  output        io_port_out_valid,
  output [15:0] io_port_out_bits,
  output [15:0] io_to_cell_bits
);
  reg  reg_0_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_0;
  reg [15:0] reg_0_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_1;
  reg  reg_1_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_2;
  reg [15:0] reg_1_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_3;
  reg  reg_2_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_4;
  reg [15:0] reg_2_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_5;
  reg  reg_3_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_6;
  reg [15:0] reg_3_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_7;
  reg  reg_4_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_8;
  reg [15:0] reg_4_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_9;
  reg  reg_5_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_10;
  reg [15:0] reg_5_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_11;
  reg  reg_6_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_12;
  reg [15:0] reg_6_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_13;
  reg  reg_7_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_14;
  reg [15:0] reg_7_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_15;
  reg  reg_8_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_16;
  reg [15:0] reg_8_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_17;
  reg  reg_9_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_18;
  reg [15:0] reg_9_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_19;
  reg  reg_10_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_20;
  reg [15:0] reg_10_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_21;
  reg  reg_11_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_22;
  reg [15:0] reg_11_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_23;
  reg [15:0] to_cell_delay1_bits; // @[pe_modules.scala 83:31]
  reg [31:0] _RAND_24;
  reg [15:0] to_cell_delay2_bits; // @[pe_modules.scala 84:31]
  reg [31:0] _RAND_25;
  assign io_port_out_valid = reg_11_valid; // @[pe_modules.scala 91:15]
  assign io_port_out_bits = reg_11_bits; // @[pe_modules.scala 91:15]
  assign io_to_cell_bits = to_cell_delay2_bits; // @[pe_modules.scala 92:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_0_bits = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_1_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_1_bits = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_2_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_2_bits = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_3_valid = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_3_bits = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_4_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_4_bits = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_5_valid = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_5_bits = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_6_valid = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_6_bits = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  reg_7_valid = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  reg_7_bits = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  reg_8_valid = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  reg_8_bits = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  reg_9_valid = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  reg_9_bits = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  reg_10_valid = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  reg_10_bits = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  reg_11_valid = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  reg_11_bits = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  to_cell_delay1_bits = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  to_cell_delay2_bits = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_0_valid <= 1'h0;
    end else begin
      reg_0_valid <= io_port_in_valid;
    end
    if (reset) begin
      reg_0_bits <= 16'h0;
    end else begin
      reg_0_bits <= io_port_in_bits;
    end
    if (reset) begin
      reg_1_valid <= 1'h0;
    end else begin
      reg_1_valid <= reg_0_valid;
    end
    if (reset) begin
      reg_1_bits <= 16'h0;
    end else begin
      reg_1_bits <= reg_0_bits;
    end
    if (reset) begin
      reg_2_valid <= 1'h0;
    end else begin
      reg_2_valid <= reg_1_valid;
    end
    if (reset) begin
      reg_2_bits <= 16'h0;
    end else begin
      reg_2_bits <= reg_1_bits;
    end
    if (reset) begin
      reg_3_valid <= 1'h0;
    end else begin
      reg_3_valid <= reg_2_valid;
    end
    if (reset) begin
      reg_3_bits <= 16'h0;
    end else begin
      reg_3_bits <= reg_2_bits;
    end
    if (reset) begin
      reg_4_valid <= 1'h0;
    end else begin
      reg_4_valid <= reg_3_valid;
    end
    if (reset) begin
      reg_4_bits <= 16'h0;
    end else begin
      reg_4_bits <= reg_3_bits;
    end
    if (reset) begin
      reg_5_valid <= 1'h0;
    end else begin
      reg_5_valid <= reg_4_valid;
    end
    if (reset) begin
      reg_5_bits <= 16'h0;
    end else begin
      reg_5_bits <= reg_4_bits;
    end
    if (reset) begin
      reg_6_valid <= 1'h0;
    end else begin
      reg_6_valid <= reg_5_valid;
    end
    if (reset) begin
      reg_6_bits <= 16'h0;
    end else begin
      reg_6_bits <= reg_5_bits;
    end
    if (reset) begin
      reg_7_valid <= 1'h0;
    end else begin
      reg_7_valid <= reg_6_valid;
    end
    if (reset) begin
      reg_7_bits <= 16'h0;
    end else begin
      reg_7_bits <= reg_6_bits;
    end
    if (reset) begin
      reg_8_valid <= 1'h0;
    end else begin
      reg_8_valid <= reg_7_valid;
    end
    if (reset) begin
      reg_8_bits <= 16'h0;
    end else begin
      reg_8_bits <= reg_7_bits;
    end
    if (reset) begin
      reg_9_valid <= 1'h0;
    end else begin
      reg_9_valid <= reg_8_valid;
    end
    if (reset) begin
      reg_9_bits <= 16'h0;
    end else begin
      reg_9_bits <= reg_8_bits;
    end
    if (reset) begin
      reg_10_valid <= 1'h0;
    end else begin
      reg_10_valid <= reg_9_valid;
    end
    if (reset) begin
      reg_10_bits <= 16'h0;
    end else begin
      reg_10_bits <= reg_9_bits;
    end
    if (reset) begin
      reg_11_valid <= 1'h0;
    end else begin
      reg_11_valid <= reg_10_valid;
    end
    if (reset) begin
      reg_11_bits <= 16'h0;
    end else begin
      reg_11_bits <= reg_10_bits;
    end
    if (reset) begin
      to_cell_delay1_bits <= 16'h0;
    end else begin
      to_cell_delay1_bits <= reg_0_bits;
    end
    if (reset) begin
      to_cell_delay2_bits <= 16'h0;
    end else begin
      to_cell_delay2_bits <= to_cell_delay1_bits;
    end
  end
endmodule
module PE(
  input         clock,
  input         reset,
  input         io_data_2_in_valid,
  input  [15:0] io_data_2_in_bits,
  output        io_data_2_out_valid,
  output [15:0] io_data_2_out_bits,
  input         io_data_1_in_valid,
  input  [15:0] io_data_1_in_bits,
  output        io_data_1_out_valid,
  output [15:0] io_data_1_out_bits,
  input         io_data_0_in_valid,
  input  [15:0] io_data_0_in_bits,
  output        io_data_0_out_valid,
  output [15:0] io_data_0_out_bits,
  input         io_sig_stat2trans
);
  wire  ComputeCell_Latency_clock; // @[pe.scala 37:104]
  wire  ComputeCell_Latency_reset; // @[pe.scala 37:104]
  wire [15:0] ComputeCell_Latency_io_data_2_in; // @[pe.scala 37:104]
  wire [15:0] ComputeCell_Latency_io_data_1_in; // @[pe.scala 37:104]
  wire [15:0] ComputeCell_Latency_io_data_0_in; // @[pe.scala 37:104]
  wire [15:0] ComputeCell_Latency_io_data_0_out; // @[pe.scala 37:104]
  wire  SystolicOutput_io_port_in_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_port_in_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_port_out_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_port_out_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_from_cell_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_from_cell_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_to_cell_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_to_cell_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_clock; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_reset; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_port_in_valid; // @[pe.scala 39:11]
  wire [15:0] StationaryInput_Pipeline_io_port_in_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_port_out_valid; // @[pe.scala 39:11]
  wire [15:0] StationaryInput_Pipeline_io_port_out_bits; // @[pe.scala 39:11]
  wire [15:0] StationaryInput_Pipeline_io_to_cell_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_sig_stat2trans; // @[pe.scala 39:11]
  wire  SystolicInput_clock; // @[pe.scala 39:11]
  wire  SystolicInput_reset; // @[pe.scala 39:11]
  wire  SystolicInput_io_port_in_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicInput_io_port_in_bits; // @[pe.scala 39:11]
  wire  SystolicInput_io_port_out_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicInput_io_port_out_bits; // @[pe.scala 39:11]
  wire [15:0] SystolicInput_io_to_cell_bits; // @[pe.scala 39:11]
  reg  _T_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  _T_4; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  _T_5; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  _T_6; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  _T_7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  _T_8; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  _T_9; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  _T_10; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  _T_11; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  _T_12; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg  _T_13; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  _T_14; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  ComputeCell_Latency ComputeCell_Latency ( // @[pe.scala 37:104]
    .clock(ComputeCell_Latency_clock),
    .reset(ComputeCell_Latency_reset),
    .io_data_2_in(ComputeCell_Latency_io_data_2_in),
    .io_data_1_in(ComputeCell_Latency_io_data_1_in),
    .io_data_0_in(ComputeCell_Latency_io_data_0_in),
    .io_data_0_out(ComputeCell_Latency_io_data_0_out)
  );
  SystolicOutput SystolicOutput ( // @[pe.scala 39:11]
    .io_port_in_valid(SystolicOutput_io_port_in_valid),
    .io_port_in_bits(SystolicOutput_io_port_in_bits),
    .io_port_out_valid(SystolicOutput_io_port_out_valid),
    .io_port_out_bits(SystolicOutput_io_port_out_bits),
    .io_from_cell_valid(SystolicOutput_io_from_cell_valid),
    .io_from_cell_bits(SystolicOutput_io_from_cell_bits),
    .io_to_cell_valid(SystolicOutput_io_to_cell_valid),
    .io_to_cell_bits(SystolicOutput_io_to_cell_bits)
  );
  StationaryInput_Pipeline StationaryInput_Pipeline ( // @[pe.scala 39:11]
    .clock(StationaryInput_Pipeline_clock),
    .reset(StationaryInput_Pipeline_reset),
    .io_port_in_valid(StationaryInput_Pipeline_io_port_in_valid),
    .io_port_in_bits(StationaryInput_Pipeline_io_port_in_bits),
    .io_port_out_valid(StationaryInput_Pipeline_io_port_out_valid),
    .io_port_out_bits(StationaryInput_Pipeline_io_port_out_bits),
    .io_to_cell_bits(StationaryInput_Pipeline_io_to_cell_bits),
    .io_sig_stat2trans(StationaryInput_Pipeline_io_sig_stat2trans)
  );
  SystolicInput SystolicInput ( // @[pe.scala 39:11]
    .clock(SystolicInput_clock),
    .reset(SystolicInput_reset),
    .io_port_in_valid(SystolicInput_io_port_in_valid),
    .io_port_in_bits(SystolicInput_io_port_in_bits),
    .io_port_out_valid(SystolicInput_io_port_out_valid),
    .io_port_out_bits(SystolicInput_io_port_out_bits),
    .io_to_cell_bits(SystolicInput_io_to_cell_bits)
  );
  assign io_data_2_out_valid = SystolicInput_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_2_out_bits = SystolicInput_io_port_out_bits; // @[pe.scala 42:17]
  assign io_data_1_out_valid = StationaryInput_Pipeline_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_1_out_bits = StationaryInput_Pipeline_io_port_out_bits; // @[pe.scala 42:17]
  assign io_data_0_out_valid = SystolicOutput_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_0_out_bits = SystolicOutput_io_port_out_bits; // @[pe.scala 42:17]
  assign ComputeCell_Latency_clock = clock;
  assign ComputeCell_Latency_reset = reset;
  assign ComputeCell_Latency_io_data_2_in = SystolicInput_io_to_cell_bits; // @[pe.scala 43:19]
  assign ComputeCell_Latency_io_data_1_in = StationaryInput_Pipeline_io_to_cell_bits; // @[pe.scala 43:19]
  assign ComputeCell_Latency_io_data_0_in = SystolicOutput_io_to_cell_bits; // @[pe.scala 43:19]
  assign SystolicOutput_io_port_in_valid = io_data_0_in_valid; // @[pe.scala 42:17]
  assign SystolicOutput_io_port_in_bits = io_data_0_in_bits; // @[pe.scala 42:17]
  assign SystolicOutput_io_from_cell_valid = _T_14; // @[pe.scala 46:34]
  assign SystolicOutput_io_from_cell_bits = ComputeCell_Latency_io_data_0_out; // @[pe.scala 45:33]
  assign StationaryInput_Pipeline_clock = clock;
  assign StationaryInput_Pipeline_reset = reset;
  assign StationaryInput_Pipeline_io_port_in_valid = io_data_1_in_valid; // @[pe.scala 42:17]
  assign StationaryInput_Pipeline_io_port_in_bits = io_data_1_in_bits; // @[pe.scala 42:17]
  assign StationaryInput_Pipeline_io_sig_stat2trans = io_sig_stat2trans; // @[pe.scala 50:33]
  assign SystolicInput_clock = clock;
  assign SystolicInput_reset = reset;
  assign SystolicInput_io_port_in_valid = io_data_2_in_valid; // @[pe.scala 42:17]
  assign SystolicInput_io_port_in_bits = io_data_2_in_bits; // @[pe.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_5 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_6 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_7 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_8 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_9 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_10 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_11 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_12 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_13 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_14 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_3 <= SystolicOutput_io_to_cell_valid;
    _T_4 <= _T_3;
    _T_5 <= _T_4;
    _T_6 <= _T_5;
    _T_7 <= _T_6;
    _T_8 <= _T_7;
    _T_9 <= _T_8;
    _T_10 <= _T_9;
    _T_11 <= _T_10;
    _T_12 <= _T_11;
    _T_13 <= _T_12;
    _T_14 <= _T_13;
  end
endmodule
module PENetwork(
  input         io_to_pes_0_out_valid,
  input  [15:0] io_to_pes_0_out_bits,
  output        io_to_pes_1_in_valid,
  output [15:0] io_to_pes_1_in_bits,
  input         io_to_pes_1_out_valid,
  input  [15:0] io_to_pes_1_out_bits,
  output        io_to_pes_2_in_valid,
  output [15:0] io_to_pes_2_in_bits,
  input         io_to_pes_2_out_valid,
  input  [15:0] io_to_pes_2_out_bits,
  output        io_to_pes_3_in_valid,
  output [15:0] io_to_pes_3_in_bits,
  input         io_to_pes_3_out_valid,
  input  [15:0] io_to_pes_3_out_bits,
  output        io_to_pes_4_in_valid,
  output [15:0] io_to_pes_4_in_bits,
  input         io_to_pes_4_out_valid,
  input  [15:0] io_to_pes_4_out_bits,
  output        io_to_pes_5_in_valid,
  output [15:0] io_to_pes_5_in_bits,
  input         io_to_pes_5_out_valid,
  input  [15:0] io_to_pes_5_out_bits,
  output        io_to_pes_6_in_valid,
  output [15:0] io_to_pes_6_in_bits,
  input         io_to_pes_6_out_valid,
  input  [15:0] io_to_pes_6_out_bits,
  output        io_to_pes_7_in_valid,
  output [15:0] io_to_pes_7_in_bits,
  input         io_to_pes_7_out_valid,
  input  [15:0] io_to_pes_7_out_bits,
  output        io_to_pes_8_in_valid,
  output [15:0] io_to_pes_8_in_bits,
  input         io_to_pes_8_out_valid,
  input  [15:0] io_to_pes_8_out_bits,
  output        io_to_pes_9_in_valid,
  output [15:0] io_to_pes_9_in_bits,
  input         io_to_pes_9_out_valid,
  input  [15:0] io_to_pes_9_out_bits,
  output        io_to_pes_10_in_valid,
  output [15:0] io_to_pes_10_in_bits,
  input         io_to_pes_10_out_valid,
  input  [15:0] io_to_pes_10_out_bits,
  output        io_to_pes_11_in_valid,
  output [15:0] io_to_pes_11_in_bits,
  input         io_to_pes_11_out_valid,
  input  [15:0] io_to_pes_11_out_bits,
  output        io_to_pes_12_in_valid,
  output [15:0] io_to_pes_12_in_bits,
  input         io_to_pes_12_out_valid,
  input  [15:0] io_to_pes_12_out_bits,
  output        io_to_pes_13_in_valid,
  output [15:0] io_to_pes_13_in_bits,
  input         io_to_pes_13_out_valid,
  input  [15:0] io_to_pes_13_out_bits,
  output        io_to_pes_14_in_valid,
  output [15:0] io_to_pes_14_in_bits,
  input         io_to_pes_14_out_valid,
  input  [15:0] io_to_pes_14_out_bits,
  output        io_to_pes_15_in_valid,
  output [15:0] io_to_pes_15_in_bits,
  input         io_to_pes_15_out_valid,
  input  [15:0] io_to_pes_15_out_bits,
  output        io_to_mem_valid,
  output [15:0] io_to_mem_bits
);
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_8_in_valid = io_to_pes_7_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_9_in_valid = io_to_pes_8_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_10_in_valid = io_to_pes_9_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_11_in_valid = io_to_pes_10_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_11_in_bits = io_to_pes_10_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_12_in_valid = io_to_pes_11_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_12_in_bits = io_to_pes_11_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_13_in_valid = io_to_pes_12_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_13_in_bits = io_to_pes_12_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_14_in_valid = io_to_pes_13_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_14_in_bits = io_to_pes_13_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_15_in_valid = io_to_pes_14_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_15_in_bits = io_to_pes_14_out_bits; // @[pearray.scala 38:23]
  assign io_to_mem_valid = io_to_pes_15_out_valid; // @[pearray.scala 45:17]
  assign io_to_mem_bits = io_to_pes_15_out_bits; // @[pearray.scala 45:17]
endmodule
module PENetwork_16(
  output        io_to_pes_0_in_valid,
  output [15:0] io_to_pes_0_in_bits,
  input         io_to_pes_0_out_valid,
  input  [15:0] io_to_pes_0_out_bits,
  output        io_to_pes_1_in_valid,
  output [15:0] io_to_pes_1_in_bits,
  input         io_to_pes_1_out_valid,
  input  [15:0] io_to_pes_1_out_bits,
  output        io_to_pes_2_in_valid,
  output [15:0] io_to_pes_2_in_bits,
  input         io_to_pes_2_out_valid,
  input  [15:0] io_to_pes_2_out_bits,
  output        io_to_pes_3_in_valid,
  output [15:0] io_to_pes_3_in_bits,
  input         io_to_pes_3_out_valid,
  input  [15:0] io_to_pes_3_out_bits,
  output        io_to_pes_4_in_valid,
  output [15:0] io_to_pes_4_in_bits,
  input         io_to_pes_4_out_valid,
  input  [15:0] io_to_pes_4_out_bits,
  output        io_to_pes_5_in_valid,
  output [15:0] io_to_pes_5_in_bits,
  input         io_to_pes_5_out_valid,
  input  [15:0] io_to_pes_5_out_bits,
  output        io_to_pes_6_in_valid,
  output [15:0] io_to_pes_6_in_bits,
  input         io_to_pes_6_out_valid,
  input  [15:0] io_to_pes_6_out_bits,
  output        io_to_pes_7_in_valid,
  output [15:0] io_to_pes_7_in_bits,
  input         io_to_pes_7_out_valid,
  input  [15:0] io_to_pes_7_out_bits,
  output        io_to_pes_8_in_valid,
  output [15:0] io_to_pes_8_in_bits,
  input         io_to_pes_8_out_valid,
  input  [15:0] io_to_pes_8_out_bits,
  output        io_to_pes_9_in_valid,
  output [15:0] io_to_pes_9_in_bits,
  input         io_to_pes_9_out_valid,
  input  [15:0] io_to_pes_9_out_bits,
  output        io_to_pes_10_in_valid,
  output [15:0] io_to_pes_10_in_bits,
  input         io_to_pes_10_out_valid,
  input  [15:0] io_to_pes_10_out_bits,
  output        io_to_pes_11_in_valid,
  output [15:0] io_to_pes_11_in_bits,
  input         io_to_pes_11_out_valid,
  input  [15:0] io_to_pes_11_out_bits,
  output        io_to_pes_12_in_valid,
  output [15:0] io_to_pes_12_in_bits,
  input         io_to_pes_12_out_valid,
  input  [15:0] io_to_pes_12_out_bits,
  output        io_to_pes_13_in_valid,
  output [15:0] io_to_pes_13_in_bits,
  input         io_to_pes_13_out_valid,
  input  [15:0] io_to_pes_13_out_bits,
  output        io_to_pes_14_in_valid,
  output [15:0] io_to_pes_14_in_bits,
  input         io_to_pes_14_out_valid,
  input  [15:0] io_to_pes_14_out_bits,
  output        io_to_pes_15_in_valid,
  output [15:0] io_to_pes_15_in_bits,
  input         io_to_mem_valid,
  input  [15:0] io_to_mem_bits
);
  assign io_to_pes_0_in_valid = io_to_mem_valid; // @[pearray.scala 41:23]
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pearray.scala 41:23]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_8_in_valid = io_to_pes_7_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_9_in_valid = io_to_pes_8_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_10_in_valid = io_to_pes_9_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_11_in_valid = io_to_pes_10_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_11_in_bits = io_to_pes_10_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_12_in_valid = io_to_pes_11_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_12_in_bits = io_to_pes_11_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_13_in_valid = io_to_pes_12_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_13_in_bits = io_to_pes_12_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_14_in_valid = io_to_pes_13_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_14_in_bits = io_to_pes_13_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_15_in_valid = io_to_pes_14_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_15_in_bits = io_to_pes_14_out_bits; // @[pearray.scala 38:23]
endmodule
module Reduction_Dummy(
  input  [15:0] io_in_a,
  input  [15:0] io_in_b,
  output [15:0] io_out
);
  assign io_out = io_in_a + io_in_b; // @[cell.scala 275:10]
endmodule
module MultiDimMem(
  input         clock,
  input         reset,
  input         io_rd_addr_valid,
  input  [1:0]  io_rd_addr_bits_0,
  input  [1:0]  io_rd_addr_bits_1,
  input  [1:0]  io_rd_addr_bits_2,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input         io_wr_addr_valid,
  input  [1:0]  io_wr_addr_bits_0,
  input  [1:0]  io_wr_addr_bits_1,
  input  [1:0]  io_wr_addr_bits_2,
  input  [1:0]  io_wr_addr_bits_3,
  input  [1:0]  io_wr_addr_bits_4,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits,
  input         io_wr_update
);
  reg [16:0] mem [0:1439]; // @[mem.scala 131:24]
  reg [31:0] _RAND_0;
  wire [16:0] mem_mem_output_data; // @[mem.scala 131:24]
  wire [10:0] mem_mem_output_addr; // @[mem.scala 131:24]
  reg [31:0] _RAND_1;
  wire [16:0] mem__T_79_data; // @[mem.scala 131:24]
  wire [10:0] mem__T_79_addr; // @[mem.scala 131:24]
  wire  mem__T_79_mask; // @[mem.scala 131:24]
  wire  mem__T_79_en; // @[mem.scala 131:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [10:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [15:0] Reduction_Dummy_io_in_a; // @[mem.scala 183:30]
  wire [15:0] Reduction_Dummy_io_in_b; // @[mem.scala 183:30]
  wire [15:0] Reduction_Dummy_io_out; // @[mem.scala 183:30]
  reg  rd_addr_reg_valid; // @[mem.scala 132:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 132:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 132:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 132:28]
  reg [31:0] _RAND_7;
  wire [15:0] _T_8 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 143:102]
  wire  _T_9 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_11 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_13 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 143:102]
  wire  _T_14 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_16 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_18 = rd_addr_reg_bits_2 + 16'hf0; // @[mem.scala 143:102]
  wire  _T_19 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_21 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_23 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 146:46]
  wire [15:0] mem_rd_addr = _T_23 + rd_addr_reg_bits_2; // @[mem.scala 146:46]
  reg  mem_req_valid; // @[mem.scala 151:30]
  reg [31:0] _RAND_8;
  reg  wr_addr_reg_valid; // @[mem.scala 152:28]
  reg [31:0] _RAND_9;
  reg [15:0] wr_addr_reg_bits_4; // @[mem.scala 152:28]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_3; // @[mem.scala 152:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 152:28]
  reg [31:0] _RAND_12;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 152:28]
  reg [31:0] _RAND_13;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 152:28]
  reg [31:0] _RAND_14;
  wire [15:0] _T_37 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 164:102]
  wire  _T_38 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_40 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_42 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 164:102]
  wire  _T_43 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_45 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [16:0] _T_46 = {{1'd0}, wr_addr_reg_bits_2}; // @[mem.scala 164:102]
  wire  _T_48 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_50 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire [16:0] _T_51 = {{1'd0}, wr_addr_reg_bits_3}; // @[mem.scala 164:102]
  wire  _T_53 = 2'h1 == io_wr_addr_bits_3; // @[Mux.scala 68:19]
  wire  _T_55 = 2'h0 == io_wr_addr_bits_3; // @[Mux.scala 68:19]
  wire [15:0] _T_57 = wr_addr_reg_bits_4 + 16'h5a0; // @[mem.scala 164:102]
  wire  _T_58 = 2'h1 == io_wr_addr_bits_4; // @[Mux.scala 68:19]
  wire  _T_60 = 2'h0 == io_wr_addr_bits_4; // @[Mux.scala 68:19]
  wire [15:0] _T_62 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 166:46]
  wire [15:0] _T_64 = _T_62 + wr_addr_reg_bits_2; // @[mem.scala 166:46]
  wire [15:0] _T_66 = _T_64 + wr_addr_reg_bits_3; // @[mem.scala 166:46]
  wire [15:0] mem_wr_addr = _T_66 + wr_addr_reg_bits_4; // @[mem.scala 166:46]
  reg  wr_data_1_valid; // @[mem.scala 171:26]
  reg [31:0] _RAND_15;
  reg [15:0] wr_data_1_bits; // @[mem.scala 171:26]
  reg [31:0] _RAND_16;
  reg  wr_update_1; // @[mem.scala 172:28]
  reg [31:0] _RAND_17;
  wire [15:0] final_rd_addr = wr_update_1 ? mem_wr_addr : mem_rd_addr; // @[mem.scala 175:26]
  reg  wr_data_2_valid; // @[mem.scala 178:26]
  reg [31:0] _RAND_18;
  reg [15:0] wr_data_2_bits; // @[mem.scala 178:26]
  reg [31:0] _RAND_19;
  reg  wr_update_2; // @[mem.scala 179:28]
  reg [31:0] _RAND_20;
  reg [15:0] wr_addr_2; // @[mem.scala 180:26]
  reg [31:0] _RAND_21;
  reg [15:0] wr_data_final; // @[mem.scala 186:30]
  reg [31:0] _RAND_22;
  reg [15:0] wr_addr_3; // @[mem.scala 187:26]
  reg [31:0] _RAND_23;
  reg  wr_valid_3; // @[mem.scala 188:27]
  reg [31:0] _RAND_24;
  wire [16:0] _GEN_9 = {wr_valid_3, 16'h0}; // @[mem.scala 191:38]
  wire [31:0] _T_75 = {{15'd0}, _GEN_9}; // @[mem.scala 191:38]
  wire [31:0] _GEN_10 = {{16'd0}, wr_data_final}; // @[mem.scala 191:52]
  wire [31:0] _T_76 = _T_75 | _GEN_10; // @[mem.scala 191:52]
  reg  _T_82; // @[mem.scala 194:30]
  reg [31:0] _RAND_25;
  reg [15:0] _T_85; // @[mem.scala 195:29]
  reg [31:0] _RAND_26;
  Reduction_Dummy Reduction_Dummy ( // @[mem.scala 183:30]
    .io_in_a(Reduction_Dummy_io_in_a),
    .io_in_b(Reduction_Dummy_io_in_b),
    .io_out(Reduction_Dummy_io_out)
  );
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 131:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 11'h5a0 ? _RAND_1[16:0] : mem[mem_mem_output_addr]; // @[mem.scala 131:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_79_data = _T_76[16:0];
  assign mem__T_79_addr = wr_addr_3[10:0];
  assign mem__T_79_mask = 1'h1;
  assign mem__T_79_en = wr_valid_3;
  assign io_rd_data_valid = _T_82; // @[mem.scala 194:20]
  assign io_rd_data_bits = _T_85; // @[mem.scala 195:19]
  assign Reduction_Dummy_io_in_a = mem_mem_output_data[15:0]; // @[mem.scala 184:23]
  assign Reduction_Dummy_io_in_b = wr_data_2_bits; // @[mem.scala 185:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1440; initvar = initvar+1)
    mem[initvar] = _RAND_0[16:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_req_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_addr_reg_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_addr_reg_bits_4 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_3 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wr_data_1_valid = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wr_data_1_bits = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  wr_update_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wr_data_2_valid = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  wr_data_2_bits = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  wr_update_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  wr_addr_2 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  wr_data_final = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  wr_addr_3 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  wr_valid_3 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_82 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_85 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_79_en & mem__T_79_mask) begin
      mem[mem__T_79_addr] <= mem__T_79_data; // @[mem.scala 131:24]
    end
    if (wr_update_1) begin
      mem_mem_output_en_pipe_0 <= wr_addr_reg_valid;
    end else begin
      mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    end
    if (wr_update_1 ? wr_addr_reg_valid : rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= final_rd_addr[10:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_21) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_19) begin
      rd_addr_reg_bits_2 <= _T_18;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_16) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= _T_13;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_11) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= _T_8;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_valid <= 1'h0;
    end else begin
      wr_addr_reg_valid <= io_wr_addr_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_4 <= 16'h0;
    end else if (_T_60) begin
      wr_addr_reg_bits_4 <= 16'h0;
    end else if (_T_58) begin
      wr_addr_reg_bits_4 <= _T_57;
    end
    if (reset) begin
      wr_addr_reg_bits_3 <= 16'h0;
    end else if (_T_55) begin
      wr_addr_reg_bits_3 <= 16'h0;
    end else if (_T_53) begin
      wr_addr_reg_bits_3 <= _T_51[15:0];
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_50) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_48) begin
      wr_addr_reg_bits_2 <= _T_46[15:0];
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_45) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_43) begin
      wr_addr_reg_bits_1 <= _T_42;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_40) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_38) begin
      wr_addr_reg_bits_0 <= _T_37;
    end
    if (reset) begin
      wr_data_1_valid <= 1'h0;
    end else begin
      wr_data_1_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_1_bits <= 16'h0;
    end else begin
      wr_data_1_bits <= io_wr_data_bits;
    end
    if (reset) begin
      wr_update_1 <= 1'h0;
    end else begin
      wr_update_1 <= io_wr_update;
    end
    if (reset) begin
      wr_data_2_valid <= 1'h0;
    end else begin
      wr_data_2_valid <= wr_data_1_valid;
    end
    if (reset) begin
      wr_data_2_bits <= 16'h0;
    end else begin
      wr_data_2_bits <= wr_data_1_bits;
    end
    if (reset) begin
      wr_update_2 <= 1'h0;
    end else begin
      wr_update_2 <= wr_update_1;
    end
    if (reset) begin
      wr_addr_2 <= 16'h0;
    end else begin
      wr_addr_2 <= mem_wr_addr;
    end
    if (wr_update_2) begin
      wr_data_final <= Reduction_Dummy_io_out;
    end else begin
      wr_data_final <= wr_data_2_bits;
    end
    if (reset) begin
      wr_addr_3 <= 16'h0;
    end else begin
      wr_addr_3 <= wr_addr_2;
    end
    wr_valid_3 <= wr_data_2_valid;
    _T_82 <= mem_req_valid & mem_mem_output_data[16];
    if (mem_req_valid) begin
      _T_85 <= mem_mem_output_data[15:0];
    end else begin
      _T_85 <= 16'h0;
    end
  end
endmodule
module MultiDimTime_5(
  input        clock,
  input        reset,
  input        io_in,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2
);
  reg [15:0] regs_0; // @[mem.scala 81:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 81:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 81:12]
  reg [31:0] _RAND_2;
  wire [15:0] _GEN_6 = {{15'd0}, io_in}; // @[mem.scala 95:42]
  wire [15:0] _T_1 = regs_0 + _GEN_6; // @[mem.scala 95:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 95:48]
  wire [15:0] _T_3 = regs_1 + _GEN_6; // @[mem.scala 95:42]
  wire  back_1 = _T_3 == 16'h14; // @[mem.scala 95:48]
  wire [15:0] _T_5 = regs_2 + _GEN_6; // @[mem.scala 95:42]
  wire  back_2 = _T_5 == 16'h6; // @[mem.scala 95:48]
  wire  _T_6 = ~back_0; // @[mem.scala 102:20]
  wire [1:0] _T_7 = {_T_6, 1'h0}; // @[mem.scala 102:31]
  wire  _T_8 = ~back_1; // @[mem.scala 102:40]
  wire [1:0] _GEN_9 = {{1'd0}, _T_8}; // @[mem.scala 102:37]
  wire  _T_12 = back_0 & back_1; // @[mem.scala 101:46]
  wire  _T_13 = ~_T_12; // @[mem.scala 102:20]
  wire [1:0] _T_14 = {_T_13, 1'h0}; // @[mem.scala 102:31]
  wire  _T_15 = ~back_2; // @[mem.scala 102:40]
  wire [1:0] _GEN_11 = {{1'd0}, _T_15}; // @[mem.scala 102:37]
  wire  _GEN_5 = back_0 ? 1'h0 : io_in; // @[mem.scala 112:16]
  assign io_out_0 = {{1'd0}, _GEN_5}; // @[mem.scala 114:15 mem.scala 117:15]
  assign io_out_1 = _T_7 | _GEN_9; // @[mem.scala 102:15]
  assign io_out_2 = _T_14 | _GEN_11; // @[mem.scala 102:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (_T_12) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
  end
endmodule
module MemController(
  input         clock,
  input         reset,
  input         io_rd_valid,
  input         io_wr_valid,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 33:19]
  wire  MultiDimMem_reset; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 33:19]
  wire [15:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 33:19]
  wire  MultiDimMem_io_wr_addr_valid; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_3; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_4; // @[mem.scala 33:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 33:19]
  wire [15:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 33:19]
  wire  MultiDimMem_io_wr_update; // @[mem.scala 33:19]
  wire  MultiDimTime_clock; // @[mem.scala 34:23]
  wire  MultiDimTime_reset; // @[mem.scala 34:23]
  wire  MultiDimTime_io_in; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_3; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_4; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_io_index_0; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_io_index_1; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_io_index_2; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_io_index_3; // @[mem.scala 34:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 35:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 35:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 35:23]
  wire [17:0] _T__0 = MultiDimTime_io_index_2; // @[mem.scala 63:48 mem.scala 63:48]
  wire  _T_1 = _T__0 == 18'h0; // @[mem.scala 63:79]
  wire [17:0] _T__1 = MultiDimTime_io_index_3; // @[mem.scala 63:48 mem.scala 63:48]
  wire  _T_2 = _T__1 == 18'h0; // @[mem.scala 63:79]
  wire  _T_4 = _T_1 & _T_2; // @[mem.scala 63:66]
  MultiDimMem MultiDimMem ( // @[mem.scala 33:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_valid(MultiDimMem_io_wr_addr_valid),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_addr_bits_3(MultiDimMem_io_wr_addr_bits_3),
    .io_wr_addr_bits_4(MultiDimMem_io_wr_addr_bits_4),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits),
    .io_wr_update(MultiDimMem_io_wr_update)
  );
  MultiDimTime MultiDimTime ( // @[mem.scala 34:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_out_3(MultiDimTime_io_out_3),
    .io_out_4(MultiDimTime_io_out_4),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2),
    .io_index_3(MultiDimTime_io_index_3)
  );
  MultiDimTime_5 MultiDimTime_1 ( // @[mem.scala 35:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 53:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 53:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 50:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 49:20]
  assign MultiDimMem_io_wr_addr_valid = io_wr_valid; // @[mem.scala 46:21]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_3 = MultiDimTime_io_out_3; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_4 = MultiDimTime_io_out_4; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 54:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 54:15]
  assign MultiDimMem_io_wr_update = ~_T_4; // @[mem.scala 47:17 mem.scala 63:19]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 44:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 48:14]
endmodule
module MultiDimMem_16(
  input         clock,
  input         reset,
  input         io_rd_addr_valid,
  input  [1:0]  io_rd_addr_bits_0,
  input  [1:0]  io_rd_addr_bits_1,
  input  [1:0]  io_rd_addr_bits_2,
  input  [1:0]  io_rd_addr_bits_3,
  input  [1:0]  io_rd_addr_bits_4,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input  [1:0]  io_wr_addr_bits_0,
  input  [1:0]  io_wr_addr_bits_1,
  input  [1:0]  io_wr_addr_bits_2,
  input  [1:0]  io_wr_addr_bits_3,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  reg [16:0] mem [0:1727]; // @[mem.scala 131:24]
  reg [31:0] _RAND_0;
  wire [16:0] mem_mem_output_data; // @[mem.scala 131:24]
  wire [10:0] mem_mem_output_addr; // @[mem.scala 131:24]
  reg [31:0] _RAND_1;
  wire [16:0] mem__T_88_data; // @[mem.scala 131:24]
  wire [10:0] mem__T_88_addr; // @[mem.scala 131:24]
  wire  mem__T_88_mask; // @[mem.scala 131:24]
  wire  mem__T_88_en; // @[mem.scala 131:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [10:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [15:0] Reduction_Dummy_io_in_a; // @[mem.scala 183:30]
  wire [15:0] Reduction_Dummy_io_in_b; // @[mem.scala 183:30]
  wire [15:0] Reduction_Dummy_io_out; // @[mem.scala 183:30]
  reg  rd_addr_reg_valid; // @[mem.scala 132:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_4; // @[mem.scala 132:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_3; // @[mem.scala 132:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 132:28]
  reg [31:0] _RAND_7;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 132:28]
  reg [31:0] _RAND_8;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 132:28]
  reg [31:0] _RAND_9;
  wire [15:0] _T_12 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 143:102]
  wire  _T_13 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_15 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_17 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 143:102]
  wire  _T_18 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_20 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_22 = rd_addr_reg_bits_2 + 16'hc0; // @[mem.scala 143:102]
  wire  _T_23 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_25 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_27 = rd_addr_reg_bits_3 + 16'h240; // @[mem.scala 143:102]
  wire  _T_28 = 2'h1 == io_rd_addr_bits_3; // @[Mux.scala 68:19]
  wire  _T_30 = 2'h0 == io_rd_addr_bits_3; // @[Mux.scala 68:19]
  wire [16:0] _T_31 = {{1'd0}, rd_addr_reg_bits_4}; // @[mem.scala 143:102]
  wire  _T_33 = 2'h1 == io_rd_addr_bits_4; // @[Mux.scala 68:19]
  wire  _T_35 = 2'h0 == io_rd_addr_bits_4; // @[Mux.scala 68:19]
  wire [15:0] _T_37 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 146:46]
  wire [15:0] _T_39 = _T_37 + rd_addr_reg_bits_2; // @[mem.scala 146:46]
  wire [15:0] _T_41 = _T_39 + rd_addr_reg_bits_3; // @[mem.scala 146:46]
  wire [15:0] mem_rd_addr = _T_41 + rd_addr_reg_bits_4; // @[mem.scala 146:46]
  reg  mem_req_valid; // @[mem.scala 151:30]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_3; // @[mem.scala 152:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 152:28]
  reg [31:0] _RAND_12;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 152:28]
  reg [31:0] _RAND_13;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 152:28]
  reg [31:0] _RAND_14;
  wire [15:0] _T_53 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 164:102]
  wire  _T_54 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_56 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_58 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 164:102]
  wire  _T_59 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_61 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_63 = wr_addr_reg_bits_2 + 16'hc0; // @[mem.scala 164:102]
  wire  _T_64 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_66 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_68 = wr_addr_reg_bits_3 + 16'h240; // @[mem.scala 164:102]
  wire  _T_69 = 2'h1 == io_wr_addr_bits_3; // @[Mux.scala 68:19]
  wire  _T_71 = 2'h0 == io_wr_addr_bits_3; // @[Mux.scala 68:19]
  wire [15:0] _T_73 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 166:46]
  wire [15:0] _T_75 = _T_73 + wr_addr_reg_bits_2; // @[mem.scala 166:46]
  wire [15:0] mem_wr_addr = _T_75 + wr_addr_reg_bits_3; // @[mem.scala 166:46]
  reg  wr_data_1_valid; // @[mem.scala 171:26]
  reg [31:0] _RAND_15;
  reg [15:0] wr_data_1_bits; // @[mem.scala 171:26]
  reg [31:0] _RAND_16;
  reg  wr_data_2_valid; // @[mem.scala 178:26]
  reg [31:0] _RAND_17;
  reg [15:0] wr_data_2_bits; // @[mem.scala 178:26]
  reg [31:0] _RAND_18;
  reg [15:0] wr_addr_2; // @[mem.scala 180:26]
  reg [31:0] _RAND_19;
  reg [15:0] wr_data_final; // @[mem.scala 186:30]
  reg [31:0] _RAND_20;
  reg [15:0] wr_addr_3; // @[mem.scala 187:26]
  reg [31:0] _RAND_21;
  reg  wr_valid_3; // @[mem.scala 188:27]
  reg [31:0] _RAND_22;
  wire [16:0] _GEN_9 = {wr_valid_3, 16'h0}; // @[mem.scala 191:38]
  wire [31:0] _T_84 = {{15'd0}, _GEN_9}; // @[mem.scala 191:38]
  wire [31:0] _GEN_10 = {{16'd0}, wr_data_final}; // @[mem.scala 191:52]
  wire [31:0] _T_85 = _T_84 | _GEN_10; // @[mem.scala 191:52]
  reg  _T_91; // @[mem.scala 194:30]
  reg [31:0] _RAND_23;
  reg [15:0] _T_94; // @[mem.scala 195:29]
  reg [31:0] _RAND_24;
  Reduction_Dummy Reduction_Dummy ( // @[mem.scala 183:30]
    .io_in_a(Reduction_Dummy_io_in_a),
    .io_in_b(Reduction_Dummy_io_in_b),
    .io_out(Reduction_Dummy_io_out)
  );
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 131:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 11'h6c0 ? _RAND_1[16:0] : mem[mem_mem_output_addr]; // @[mem.scala 131:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_88_data = _T_85[16:0];
  assign mem__T_88_addr = wr_addr_3[10:0];
  assign mem__T_88_mask = 1'h1;
  assign mem__T_88_en = wr_valid_3;
  assign io_rd_data_valid = _T_91; // @[mem.scala 194:20]
  assign io_rd_data_bits = _T_94; // @[mem.scala 195:19]
  assign Reduction_Dummy_io_in_a = mem_mem_output_data[15:0]; // @[mem.scala 184:23]
  assign Reduction_Dummy_io_in_b = wr_data_2_bits; // @[mem.scala 185:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1728; initvar = initvar+1)
    mem[initvar] = _RAND_0[16:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_4 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_3 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_req_valid = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_3 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wr_data_1_valid = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wr_data_1_bits = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  wr_data_2_valid = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wr_data_2_bits = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  wr_addr_2 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  wr_data_final = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  wr_addr_3 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  wr_valid_3 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_91 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_94 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_88_en & mem__T_88_mask) begin
      mem[mem__T_88_addr] <= mem__T_88_data; // @[mem.scala 131:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[10:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_4 <= 16'h0;
    end else if (_T_35) begin
      rd_addr_reg_bits_4 <= 16'h0;
    end else if (_T_33) begin
      rd_addr_reg_bits_4 <= _T_31[15:0];
    end
    if (reset) begin
      rd_addr_reg_bits_3 <= 16'h0;
    end else if (_T_30) begin
      rd_addr_reg_bits_3 <= 16'h0;
    end else if (_T_28) begin
      rd_addr_reg_bits_3 <= _T_27;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_25) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_23) begin
      rd_addr_reg_bits_2 <= _T_22;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_20) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_18) begin
      rd_addr_reg_bits_1 <= _T_17;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_15) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_13) begin
      rd_addr_reg_bits_0 <= _T_12;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_3 <= 16'h0;
    end else if (_T_71) begin
      wr_addr_reg_bits_3 <= 16'h0;
    end else if (_T_69) begin
      wr_addr_reg_bits_3 <= _T_68;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_66) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_64) begin
      wr_addr_reg_bits_2 <= _T_63;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_61) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_59) begin
      wr_addr_reg_bits_1 <= _T_58;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_56) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_54) begin
      wr_addr_reg_bits_0 <= _T_53;
    end
    if (reset) begin
      wr_data_1_valid <= 1'h0;
    end else begin
      wr_data_1_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_1_bits <= 16'h0;
    end else begin
      wr_data_1_bits <= io_wr_data_bits;
    end
    if (reset) begin
      wr_data_2_valid <= 1'h0;
    end else begin
      wr_data_2_valid <= wr_data_1_valid;
    end
    if (reset) begin
      wr_data_2_bits <= 16'h0;
    end else begin
      wr_data_2_bits <= wr_data_1_bits;
    end
    if (reset) begin
      wr_addr_2 <= 16'h0;
    end else begin
      wr_addr_2 <= mem_wr_addr;
    end
    wr_data_final <= wr_data_2_bits;
    if (reset) begin
      wr_addr_3 <= 16'h0;
    end else begin
      wr_addr_3 <= wr_addr_2;
    end
    wr_valid_3 <= wr_data_2_valid;
    _T_91 <= mem_req_valid & mem_mem_output_data[16];
    if (mem_req_valid) begin
      _T_94 <= mem_mem_output_data[15:0];
    end else begin
      _T_94 <= 16'h0;
    end
  end
endmodule
module MultiDimTime_36(
  input        clock,
  input        reset,
  input        io_in,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2,
  output [1:0] io_out_3
);
  reg [15:0] regs_0; // @[mem.scala 81:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 81:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 81:12]
  reg [31:0] _RAND_2;
  reg [15:0] regs_3; // @[mem.scala 81:12]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_8 = {{15'd0}, io_in}; // @[mem.scala 95:42]
  wire [15:0] _T_1 = regs_0 + _GEN_8; // @[mem.scala 95:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 95:48]
  wire [15:0] _T_3 = regs_1 + _GEN_8; // @[mem.scala 95:42]
  wire  back_1 = _T_3 == 16'h10; // @[mem.scala 95:48]
  wire [15:0] _T_5 = regs_2 + _GEN_8; // @[mem.scala 95:42]
  wire  back_2 = _T_5 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_7 = regs_3 + _GEN_8; // @[mem.scala 95:42]
  wire  back_3 = _T_7 == 16'h3; // @[mem.scala 95:48]
  wire  _T_8 = ~back_0; // @[mem.scala 102:20]
  wire [1:0] _T_9 = {_T_8, 1'h0}; // @[mem.scala 102:31]
  wire  _T_10 = ~back_1; // @[mem.scala 102:40]
  wire [1:0] _GEN_12 = {{1'd0}, _T_10}; // @[mem.scala 102:37]
  wire  _T_14 = back_0 & back_1; // @[mem.scala 101:46]
  wire  _T_15 = ~_T_14; // @[mem.scala 102:20]
  wire [1:0] _T_16 = {_T_15, 1'h0}; // @[mem.scala 102:31]
  wire  _T_17 = ~back_2; // @[mem.scala 102:40]
  wire [1:0] _GEN_14 = {{1'd0}, _T_17}; // @[mem.scala 102:37]
  wire  _T_22 = _T_14 & back_2; // @[mem.scala 101:46]
  wire  _T_23 = ~_T_22; // @[mem.scala 102:20]
  wire [1:0] _T_24 = {_T_23, 1'h0}; // @[mem.scala 102:31]
  wire  _T_25 = ~back_3; // @[mem.scala 102:40]
  wire [1:0] _GEN_16 = {{1'd0}, _T_25}; // @[mem.scala 102:37]
  wire  _GEN_7 = back_0 ? 1'h0 : io_in; // @[mem.scala 112:16]
  assign io_out_0 = {{1'd0}, _GEN_7}; // @[mem.scala 114:15 mem.scala 117:15]
  assign io_out_1 = _T_9 | _GEN_12; // @[mem.scala 102:15]
  assign io_out_2 = _T_16 | _GEN_14; // @[mem.scala 102:15]
  assign io_out_3 = _T_24 | _GEN_16; // @[mem.scala 102:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (_T_14) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
    if (reset) begin
      regs_3 <= 16'h0;
    end else if (_T_22) begin
      if (back_3) begin
        regs_3 <= 16'h0;
      end else begin
        regs_3 <= _T_7;
      end
    end
  end
endmodule
module MultiDimTime_37(
  input        clock,
  input        reset,
  input        io_in,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2,
  output [1:0] io_out_3,
  output [1:0] io_out_4
);
  reg [15:0] regs_0; // @[mem.scala 81:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 81:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 81:12]
  reg [31:0] _RAND_2;
  reg [15:0] regs_3; // @[mem.scala 81:12]
  reg [31:0] _RAND_3;
  reg [15:0] regs_4; // @[mem.scala 81:12]
  reg [31:0] _RAND_4;
  wire [15:0] _GEN_10 = {{15'd0}, io_in}; // @[mem.scala 95:42]
  wire [15:0] _T_1 = regs_0 + _GEN_10; // @[mem.scala 95:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 95:48]
  wire [15:0] _T_3 = regs_1 + _GEN_10; // @[mem.scala 95:42]
  wire  back_1 = _T_3 == 16'h10; // @[mem.scala 95:48]
  wire [15:0] _T_5 = regs_2 + _GEN_10; // @[mem.scala 95:42]
  wire  back_2 = _T_5 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_7 = regs_3 + _GEN_10; // @[mem.scala 95:42]
  wire  back_3 = _T_7 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_9 = regs_4 + _GEN_10; // @[mem.scala 95:42]
  wire  back_4 = _T_9 == 16'h6; // @[mem.scala 95:48]
  wire  _T_10 = ~back_0; // @[mem.scala 102:20]
  wire [1:0] _T_11 = {_T_10, 1'h0}; // @[mem.scala 102:31]
  wire  _T_12 = ~back_1; // @[mem.scala 102:40]
  wire [1:0] _GEN_15 = {{1'd0}, _T_12}; // @[mem.scala 102:37]
  wire  _T_16 = back_0 & back_1; // @[mem.scala 101:46]
  wire  _T_17 = ~_T_16; // @[mem.scala 102:20]
  wire [1:0] _T_18 = {_T_17, 1'h0}; // @[mem.scala 102:31]
  wire  _T_19 = ~back_2; // @[mem.scala 102:40]
  wire [1:0] _GEN_17 = {{1'd0}, _T_19}; // @[mem.scala 102:37]
  wire  _T_24 = _T_16 & back_2; // @[mem.scala 101:46]
  wire  _T_25 = ~_T_24; // @[mem.scala 102:20]
  wire [1:0] _T_26 = {_T_25, 1'h0}; // @[mem.scala 102:31]
  wire  _T_27 = ~back_3; // @[mem.scala 102:40]
  wire [1:0] _GEN_19 = {{1'd0}, _T_27}; // @[mem.scala 102:37]
  wire  _T_33 = _T_24 & back_3; // @[mem.scala 101:46]
  wire  _T_34 = ~_T_33; // @[mem.scala 102:20]
  wire [1:0] _T_35 = {_T_34, 1'h0}; // @[mem.scala 102:31]
  wire  _T_36 = ~back_4; // @[mem.scala 102:40]
  wire [1:0] _GEN_21 = {{1'd0}, _T_36}; // @[mem.scala 102:37]
  wire  _GEN_9 = back_0 ? 1'h0 : io_in; // @[mem.scala 112:16]
  assign io_out_0 = {{1'd0}, _GEN_9}; // @[mem.scala 114:15 mem.scala 117:15]
  assign io_out_1 = _T_11 | _GEN_15; // @[mem.scala 102:15]
  assign io_out_2 = _T_18 | _GEN_17; // @[mem.scala 102:15]
  assign io_out_3 = _T_26 | _GEN_19; // @[mem.scala 102:15]
  assign io_out_4 = _T_35 | _GEN_21; // @[mem.scala 102:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (_T_16) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
    if (reset) begin
      regs_3 <= 16'h0;
    end else if (_T_24) begin
      if (back_3) begin
        regs_3 <= 16'h0;
      end else begin
        regs_3 <= _T_7;
      end
    end
    if (reset) begin
      regs_4 <= 16'h0;
    end else if (_T_33) begin
      if (back_4) begin
        regs_4 <= 16'h0;
      end else begin
        regs_4 <= _T_9;
      end
    end
  end
endmodule
module MemController_16(
  input         clock,
  input         reset,
  input         io_rd_valid,
  input         io_wr_valid,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 33:19]
  wire  MultiDimMem_reset; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_3; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_4; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 33:19]
  wire [15:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_3; // @[mem.scala 33:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 33:19]
  wire [15:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 33:19]
  wire  MultiDimTime_clock; // @[mem.scala 34:23]
  wire  MultiDimTime_reset; // @[mem.scala 34:23]
  wire  MultiDimTime_io_in; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_3; // @[mem.scala 34:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 35:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 35:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_3; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_4; // @[mem.scala 35:23]
  MultiDimMem_16 MultiDimMem ( // @[mem.scala 33:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_addr_bits_3(MultiDimMem_io_rd_addr_bits_3),
    .io_rd_addr_bits_4(MultiDimMem_io_rd_addr_bits_4),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_addr_bits_3(MultiDimMem_io_wr_addr_bits_3),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime_36 MultiDimTime ( // @[mem.scala 34:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_out_3(MultiDimTime_io_out_3)
  );
  MultiDimTime_37 MultiDimTime_1 ( // @[mem.scala 35:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2),
    .io_out_3(MultiDimTime_1_io_out_3),
    .io_out_4(MultiDimTime_1_io_out_4)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 53:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 53:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 50:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_3 = MultiDimTime_1_io_out_3; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_4 = MultiDimTime_1_io_out_4; // @[mem.scala 49:20]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_3 = MultiDimTime_io_out_3; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 54:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 54:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 44:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 48:14]
endmodule
module MultiDimMem_32(
  input         clock,
  input         reset,
  input         io_rd_addr_valid,
  input  [1:0]  io_rd_addr_bits_0,
  input  [1:0]  io_rd_addr_bits_1,
  input  [1:0]  io_rd_addr_bits_2,
  input  [1:0]  io_rd_addr_bits_3,
  input  [1:0]  io_rd_addr_bits_4,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input  [1:0]  io_wr_addr_bits_0,
  input  [1:0]  io_wr_addr_bits_1,
  input  [1:0]  io_wr_addr_bits_2,
  input  [1:0]  io_wr_addr_bits_3,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  reg [16:0] mem [0:6335]; // @[mem.scala 131:24]
  reg [31:0] _RAND_0;
  wire [16:0] mem_mem_output_data; // @[mem.scala 131:24]
  wire [12:0] mem_mem_output_addr; // @[mem.scala 131:24]
  reg [31:0] _RAND_1;
  wire [16:0] mem__T_88_data; // @[mem.scala 131:24]
  wire [12:0] mem__T_88_addr; // @[mem.scala 131:24]
  wire  mem__T_88_mask; // @[mem.scala 131:24]
  wire  mem__T_88_en; // @[mem.scala 131:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [12:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [15:0] Reduction_Dummy_io_in_a; // @[mem.scala 183:30]
  wire [15:0] Reduction_Dummy_io_in_b; // @[mem.scala 183:30]
  wire [15:0] Reduction_Dummy_io_out; // @[mem.scala 183:30]
  reg  rd_addr_reg_valid; // @[mem.scala 132:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_4; // @[mem.scala 132:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_3; // @[mem.scala 132:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 132:28]
  reg [31:0] _RAND_7;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 132:28]
  reg [31:0] _RAND_8;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 132:28]
  reg [31:0] _RAND_9;
  wire [15:0] _T_12 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 143:102]
  wire  _T_13 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_15 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_17 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 143:102]
  wire  _T_18 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_20 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_22 = rd_addr_reg_bits_2 + 16'h108; // @[mem.scala 143:102]
  wire  _T_23 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_25 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_27 = rd_addr_reg_bits_3 + 16'h318; // @[mem.scala 143:102]
  wire  _T_28 = 2'h1 == io_rd_addr_bits_3; // @[Mux.scala 68:19]
  wire  _T_30 = 2'h0 == io_rd_addr_bits_3; // @[Mux.scala 68:19]
  wire [15:0] _T_32 = rd_addr_reg_bits_4 + 16'h318; // @[mem.scala 143:102]
  wire  _T_33 = 2'h1 == io_rd_addr_bits_4; // @[Mux.scala 68:19]
  wire  _T_35 = 2'h0 == io_rd_addr_bits_4; // @[Mux.scala 68:19]
  wire [15:0] _T_37 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 146:46]
  wire [15:0] _T_39 = _T_37 + rd_addr_reg_bits_2; // @[mem.scala 146:46]
  wire [15:0] _T_41 = _T_39 + rd_addr_reg_bits_3; // @[mem.scala 146:46]
  wire [15:0] mem_rd_addr = _T_41 + rd_addr_reg_bits_4; // @[mem.scala 146:46]
  reg  mem_req_valid; // @[mem.scala 151:30]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_3; // @[mem.scala 152:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 152:28]
  reg [31:0] _RAND_12;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 152:28]
  reg [31:0] _RAND_13;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 152:28]
  reg [31:0] _RAND_14;
  wire [15:0] _T_53 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 164:102]
  wire  _T_54 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_56 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_58 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 164:102]
  wire  _T_59 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_61 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_63 = wr_addr_reg_bits_2 + 16'h108; // @[mem.scala 164:102]
  wire  _T_64 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_66 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_68 = wr_addr_reg_bits_3 + 16'h318; // @[mem.scala 164:102]
  wire  _T_69 = 2'h1 == io_wr_addr_bits_3; // @[Mux.scala 68:19]
  wire  _T_71 = 2'h0 == io_wr_addr_bits_3; // @[Mux.scala 68:19]
  wire [15:0] _T_73 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 166:46]
  wire [15:0] _T_75 = _T_73 + wr_addr_reg_bits_2; // @[mem.scala 166:46]
  wire [15:0] mem_wr_addr = _T_75 + wr_addr_reg_bits_3; // @[mem.scala 166:46]
  reg  wr_data_1_valid; // @[mem.scala 171:26]
  reg [31:0] _RAND_15;
  reg [15:0] wr_data_1_bits; // @[mem.scala 171:26]
  reg [31:0] _RAND_16;
  reg  wr_data_2_valid; // @[mem.scala 178:26]
  reg [31:0] _RAND_17;
  reg [15:0] wr_data_2_bits; // @[mem.scala 178:26]
  reg [31:0] _RAND_18;
  reg [15:0] wr_addr_2; // @[mem.scala 180:26]
  reg [31:0] _RAND_19;
  reg [15:0] wr_data_final; // @[mem.scala 186:30]
  reg [31:0] _RAND_20;
  reg [15:0] wr_addr_3; // @[mem.scala 187:26]
  reg [31:0] _RAND_21;
  reg  wr_valid_3; // @[mem.scala 188:27]
  reg [31:0] _RAND_22;
  wire [16:0] _GEN_9 = {wr_valid_3, 16'h0}; // @[mem.scala 191:38]
  wire [31:0] _T_84 = {{15'd0}, _GEN_9}; // @[mem.scala 191:38]
  wire [31:0] _GEN_10 = {{16'd0}, wr_data_final}; // @[mem.scala 191:52]
  wire [31:0] _T_85 = _T_84 | _GEN_10; // @[mem.scala 191:52]
  reg  _T_91; // @[mem.scala 194:30]
  reg [31:0] _RAND_23;
  reg [15:0] _T_94; // @[mem.scala 195:29]
  reg [31:0] _RAND_24;
  Reduction_Dummy Reduction_Dummy ( // @[mem.scala 183:30]
    .io_in_a(Reduction_Dummy_io_in_a),
    .io_in_b(Reduction_Dummy_io_in_b),
    .io_out(Reduction_Dummy_io_out)
  );
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 131:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 13'h18c0 ? _RAND_1[16:0] : mem[mem_mem_output_addr]; // @[mem.scala 131:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_88_data = _T_85[16:0];
  assign mem__T_88_addr = wr_addr_3[12:0];
  assign mem__T_88_mask = 1'h1;
  assign mem__T_88_en = wr_valid_3;
  assign io_rd_data_valid = _T_91; // @[mem.scala 194:20]
  assign io_rd_data_bits = _T_94; // @[mem.scala 195:19]
  assign Reduction_Dummy_io_in_a = mem_mem_output_data[15:0]; // @[mem.scala 184:23]
  assign Reduction_Dummy_io_in_b = wr_data_2_bits; // @[mem.scala 185:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 6336; initvar = initvar+1)
    mem[initvar] = _RAND_0[16:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_4 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_3 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_req_valid = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_3 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wr_data_1_valid = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wr_data_1_bits = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  wr_data_2_valid = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wr_data_2_bits = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  wr_addr_2 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  wr_data_final = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  wr_addr_3 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  wr_valid_3 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_91 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_94 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_88_en & mem__T_88_mask) begin
      mem[mem__T_88_addr] <= mem__T_88_data; // @[mem.scala 131:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[12:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_4 <= 16'h0;
    end else if (_T_35) begin
      rd_addr_reg_bits_4 <= 16'h0;
    end else if (_T_33) begin
      rd_addr_reg_bits_4 <= _T_32;
    end
    if (reset) begin
      rd_addr_reg_bits_3 <= 16'h0;
    end else if (_T_30) begin
      rd_addr_reg_bits_3 <= 16'h0;
    end else if (_T_28) begin
      rd_addr_reg_bits_3 <= _T_27;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_25) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_23) begin
      rd_addr_reg_bits_2 <= _T_22;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_20) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_18) begin
      rd_addr_reg_bits_1 <= _T_17;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_15) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_13) begin
      rd_addr_reg_bits_0 <= _T_12;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_3 <= 16'h0;
    end else if (_T_71) begin
      wr_addr_reg_bits_3 <= 16'h0;
    end else if (_T_69) begin
      wr_addr_reg_bits_3 <= _T_68;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_66) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_64) begin
      wr_addr_reg_bits_2 <= _T_63;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_61) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_59) begin
      wr_addr_reg_bits_1 <= _T_58;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_56) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_54) begin
      wr_addr_reg_bits_0 <= _T_53;
    end
    if (reset) begin
      wr_data_1_valid <= 1'h0;
    end else begin
      wr_data_1_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_1_bits <= 16'h0;
    end else begin
      wr_data_1_bits <= io_wr_data_bits;
    end
    if (reset) begin
      wr_data_2_valid <= 1'h0;
    end else begin
      wr_data_2_valid <= wr_data_1_valid;
    end
    if (reset) begin
      wr_data_2_bits <= 16'h0;
    end else begin
      wr_data_2_bits <= wr_data_1_bits;
    end
    if (reset) begin
      wr_addr_2 <= 16'h0;
    end else begin
      wr_addr_2 <= mem_wr_addr;
    end
    wr_data_final <= wr_data_2_bits;
    if (reset) begin
      wr_addr_3 <= 16'h0;
    end else begin
      wr_addr_3 <= wr_addr_2;
    end
    wr_valid_3 <= wr_data_2_valid;
    _T_91 <= mem_req_valid & mem_mem_output_data[16];
    if (mem_req_valid) begin
      _T_94 <= mem_mem_output_data[15:0];
    end else begin
      _T_94 <= 16'h0;
    end
  end
endmodule
module MultiDimTime_68(
  input        clock,
  input        reset,
  input        io_in,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2,
  output [1:0] io_out_3
);
  reg [15:0] regs_0; // @[mem.scala 81:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 81:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 81:12]
  reg [31:0] _RAND_2;
  reg [15:0] regs_3; // @[mem.scala 81:12]
  reg [31:0] _RAND_3;
  wire [15:0] _GEN_8 = {{15'd0}, io_in}; // @[mem.scala 95:42]
  wire [15:0] _T_1 = regs_0 + _GEN_8; // @[mem.scala 95:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 95:48]
  wire [15:0] _T_3 = regs_1 + _GEN_8; // @[mem.scala 95:42]
  wire  back_1 = _T_3 == 16'h16; // @[mem.scala 95:48]
  wire [15:0] _T_5 = regs_2 + _GEN_8; // @[mem.scala 95:42]
  wire  back_2 = _T_5 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_7 = regs_3 + _GEN_8; // @[mem.scala 95:42]
  wire  back_3 = _T_7 == 16'h8; // @[mem.scala 95:48]
  wire  _T_8 = ~back_0; // @[mem.scala 102:20]
  wire [1:0] _T_9 = {_T_8, 1'h0}; // @[mem.scala 102:31]
  wire  _T_10 = ~back_1; // @[mem.scala 102:40]
  wire [1:0] _GEN_12 = {{1'd0}, _T_10}; // @[mem.scala 102:37]
  wire  _T_14 = back_0 & back_1; // @[mem.scala 101:46]
  wire  _T_15 = ~_T_14; // @[mem.scala 102:20]
  wire [1:0] _T_16 = {_T_15, 1'h0}; // @[mem.scala 102:31]
  wire  _T_17 = ~back_2; // @[mem.scala 102:40]
  wire [1:0] _GEN_14 = {{1'd0}, _T_17}; // @[mem.scala 102:37]
  wire  _T_22 = _T_14 & back_2; // @[mem.scala 101:46]
  wire  _T_23 = ~_T_22; // @[mem.scala 102:20]
  wire [1:0] _T_24 = {_T_23, 1'h0}; // @[mem.scala 102:31]
  wire  _T_25 = ~back_3; // @[mem.scala 102:40]
  wire [1:0] _GEN_16 = {{1'd0}, _T_25}; // @[mem.scala 102:37]
  wire  _GEN_7 = back_0 ? 1'h0 : io_in; // @[mem.scala 112:16]
  assign io_out_0 = {{1'd0}, _GEN_7}; // @[mem.scala 114:15 mem.scala 117:15]
  assign io_out_1 = _T_9 | _GEN_12; // @[mem.scala 102:15]
  assign io_out_2 = _T_16 | _GEN_14; // @[mem.scala 102:15]
  assign io_out_3 = _T_24 | _GEN_16; // @[mem.scala 102:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (_T_14) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
    if (reset) begin
      regs_3 <= 16'h0;
    end else if (_T_22) begin
      if (back_3) begin
        regs_3 <= 16'h0;
      end else begin
        regs_3 <= _T_7;
      end
    end
  end
endmodule
module MultiDimTime_69(
  input        clock,
  input        reset,
  input        io_in,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2,
  output [1:0] io_out_3,
  output [1:0] io_out_4
);
  reg [15:0] regs_0; // @[mem.scala 81:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 81:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 81:12]
  reg [31:0] _RAND_2;
  reg [15:0] regs_3; // @[mem.scala 81:12]
  reg [31:0] _RAND_3;
  reg [15:0] regs_4; // @[mem.scala 81:12]
  reg [31:0] _RAND_4;
  wire [15:0] _GEN_10 = {{15'd0}, io_in}; // @[mem.scala 95:42]
  wire [15:0] _T_1 = regs_0 + _GEN_10; // @[mem.scala 95:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 95:48]
  wire [15:0] _T_3 = regs_1 + _GEN_10; // @[mem.scala 95:42]
  wire  back_1 = _T_3 == 16'h16; // @[mem.scala 95:48]
  wire [15:0] _T_5 = regs_2 + _GEN_10; // @[mem.scala 95:42]
  wire  back_2 = _T_5 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_7 = regs_3 + _GEN_10; // @[mem.scala 95:42]
  wire  back_3 = _T_7 == 16'h3; // @[mem.scala 95:48]
  wire [15:0] _T_9 = regs_4 + _GEN_10; // @[mem.scala 95:42]
  wire  back_4 = _T_9 == 16'h6; // @[mem.scala 95:48]
  wire  _T_10 = ~back_0; // @[mem.scala 102:20]
  wire [1:0] _T_11 = {_T_10, 1'h0}; // @[mem.scala 102:31]
  wire  _T_12 = ~back_1; // @[mem.scala 102:40]
  wire [1:0] _GEN_15 = {{1'd0}, _T_12}; // @[mem.scala 102:37]
  wire  _T_16 = back_0 & back_1; // @[mem.scala 101:46]
  wire  _T_17 = ~_T_16; // @[mem.scala 102:20]
  wire [1:0] _T_18 = {_T_17, 1'h0}; // @[mem.scala 102:31]
  wire  _T_19 = ~back_2; // @[mem.scala 102:40]
  wire [1:0] _GEN_17 = {{1'd0}, _T_19}; // @[mem.scala 102:37]
  wire  _T_24 = _T_16 & back_2; // @[mem.scala 101:46]
  wire  _T_25 = ~_T_24; // @[mem.scala 102:20]
  wire [1:0] _T_26 = {_T_25, 1'h0}; // @[mem.scala 102:31]
  wire  _T_27 = ~back_3; // @[mem.scala 102:40]
  wire [1:0] _GEN_19 = {{1'd0}, _T_27}; // @[mem.scala 102:37]
  wire  _T_33 = _T_24 & back_3; // @[mem.scala 101:46]
  wire  _T_34 = ~_T_33; // @[mem.scala 102:20]
  wire [1:0] _T_35 = {_T_34, 1'h0}; // @[mem.scala 102:31]
  wire  _T_36 = ~back_4; // @[mem.scala 102:40]
  wire [1:0] _GEN_21 = {{1'd0}, _T_36}; // @[mem.scala 102:37]
  wire  _GEN_9 = back_0 ? 1'h0 : io_in; // @[mem.scala 112:16]
  assign io_out_0 = {{1'd0}, _GEN_9}; // @[mem.scala 114:15 mem.scala 117:15]
  assign io_out_1 = _T_11 | _GEN_15; // @[mem.scala 102:15]
  assign io_out_2 = _T_18 | _GEN_17; // @[mem.scala 102:15]
  assign io_out_3 = _T_26 | _GEN_19; // @[mem.scala 102:15]
  assign io_out_4 = _T_35 | _GEN_21; // @[mem.scala 102:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (_T_16) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
    if (reset) begin
      regs_3 <= 16'h0;
    end else if (_T_24) begin
      if (back_3) begin
        regs_3 <= 16'h0;
      end else begin
        regs_3 <= _T_7;
      end
    end
    if (reset) begin
      regs_4 <= 16'h0;
    end else if (_T_33) begin
      if (back_4) begin
        regs_4 <= 16'h0;
      end else begin
        regs_4 <= _T_9;
      end
    end
  end
endmodule
module MemController_32(
  input         clock,
  input         reset,
  input         io_rd_valid,
  input         io_wr_valid,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 33:19]
  wire  MultiDimMem_reset; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_3; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_4; // @[mem.scala 33:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 33:19]
  wire [15:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 33:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_3; // @[mem.scala 33:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 33:19]
  wire [15:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 33:19]
  wire  MultiDimTime_clock; // @[mem.scala 34:23]
  wire  MultiDimTime_reset; // @[mem.scala 34:23]
  wire  MultiDimTime_io_in; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_io_out_3; // @[mem.scala 34:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 35:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 35:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_3; // @[mem.scala 35:23]
  wire [1:0] MultiDimTime_1_io_out_4; // @[mem.scala 35:23]
  MultiDimMem_32 MultiDimMem ( // @[mem.scala 33:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_addr_bits_3(MultiDimMem_io_rd_addr_bits_3),
    .io_rd_addr_bits_4(MultiDimMem_io_rd_addr_bits_4),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_addr_bits_3(MultiDimMem_io_wr_addr_bits_3),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime_68 MultiDimTime ( // @[mem.scala 34:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_out_3(MultiDimTime_io_out_3)
  );
  MultiDimTime_69 MultiDimTime_1 ( // @[mem.scala 35:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2),
    .io_out_3(MultiDimTime_1_io_out_3),
    .io_out_4(MultiDimTime_1_io_out_4)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 53:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 53:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 50:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_3 = MultiDimTime_1_io_out_3; // @[mem.scala 49:20]
  assign MultiDimMem_io_rd_addr_bits_4 = MultiDimTime_1_io_out_4; // @[mem.scala 49:20]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_addr_bits_3 = MultiDimTime_io_out_3; // @[mem.scala 45:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 54:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 54:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 44:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 48:14]
endmodule
module PEArray(
  input         clock,
  input         reset,
  input         io_data_2_in_0_valid,
  input         io_data_2_in_0_bits_valid,
  input  [15:0] io_data_2_in_0_bits_bits,
  input         io_data_2_in_1_valid,
  input         io_data_2_in_1_bits_valid,
  input  [15:0] io_data_2_in_1_bits_bits,
  input         io_data_2_in_2_valid,
  input         io_data_2_in_2_bits_valid,
  input  [15:0] io_data_2_in_2_bits_bits,
  input         io_data_2_in_3_valid,
  input         io_data_2_in_3_bits_valid,
  input  [15:0] io_data_2_in_3_bits_bits,
  input         io_data_2_in_4_valid,
  input         io_data_2_in_4_bits_valid,
  input  [15:0] io_data_2_in_4_bits_bits,
  input         io_data_2_in_5_valid,
  input         io_data_2_in_5_bits_valid,
  input  [15:0] io_data_2_in_5_bits_bits,
  input         io_data_2_in_6_valid,
  input         io_data_2_in_6_bits_valid,
  input  [15:0] io_data_2_in_6_bits_bits,
  input         io_data_2_in_7_valid,
  input         io_data_2_in_7_bits_valid,
  input  [15:0] io_data_2_in_7_bits_bits,
  input         io_data_2_in_8_valid,
  input         io_data_2_in_8_bits_valid,
  input  [15:0] io_data_2_in_8_bits_bits,
  input         io_data_2_in_9_valid,
  input         io_data_2_in_9_bits_valid,
  input  [15:0] io_data_2_in_9_bits_bits,
  input         io_data_2_in_10_valid,
  input         io_data_2_in_10_bits_valid,
  input  [15:0] io_data_2_in_10_bits_bits,
  input         io_data_2_in_11_valid,
  input         io_data_2_in_11_bits_valid,
  input  [15:0] io_data_2_in_11_bits_bits,
  input         io_data_2_in_12_valid,
  input         io_data_2_in_12_bits_valid,
  input  [15:0] io_data_2_in_12_bits_bits,
  input         io_data_2_in_13_valid,
  input         io_data_2_in_13_bits_valid,
  input  [15:0] io_data_2_in_13_bits_bits,
  input         io_data_2_in_14_valid,
  input         io_data_2_in_14_bits_valid,
  input  [15:0] io_data_2_in_14_bits_bits,
  input         io_data_2_in_15_valid,
  input         io_data_2_in_15_bits_valid,
  input  [15:0] io_data_2_in_15_bits_bits,
  input         io_data_1_in_0_valid,
  input         io_data_1_in_0_bits_valid,
  input  [15:0] io_data_1_in_0_bits_bits,
  input         io_data_1_in_1_valid,
  input         io_data_1_in_1_bits_valid,
  input  [15:0] io_data_1_in_1_bits_bits,
  input         io_data_1_in_2_valid,
  input         io_data_1_in_2_bits_valid,
  input  [15:0] io_data_1_in_2_bits_bits,
  input         io_data_1_in_3_valid,
  input         io_data_1_in_3_bits_valid,
  input  [15:0] io_data_1_in_3_bits_bits,
  input         io_data_1_in_4_valid,
  input         io_data_1_in_4_bits_valid,
  input  [15:0] io_data_1_in_4_bits_bits,
  input         io_data_1_in_5_valid,
  input         io_data_1_in_5_bits_valid,
  input  [15:0] io_data_1_in_5_bits_bits,
  input         io_data_1_in_6_valid,
  input         io_data_1_in_6_bits_valid,
  input  [15:0] io_data_1_in_6_bits_bits,
  input         io_data_1_in_7_valid,
  input         io_data_1_in_7_bits_valid,
  input  [15:0] io_data_1_in_7_bits_bits,
  input         io_data_1_in_8_valid,
  input         io_data_1_in_8_bits_valid,
  input  [15:0] io_data_1_in_8_bits_bits,
  input         io_data_1_in_9_valid,
  input         io_data_1_in_9_bits_valid,
  input  [15:0] io_data_1_in_9_bits_bits,
  input         io_data_1_in_10_valid,
  input         io_data_1_in_10_bits_valid,
  input  [15:0] io_data_1_in_10_bits_bits,
  input         io_data_1_in_11_valid,
  input         io_data_1_in_11_bits_valid,
  input  [15:0] io_data_1_in_11_bits_bits,
  input         io_data_1_in_12_valid,
  input         io_data_1_in_12_bits_valid,
  input  [15:0] io_data_1_in_12_bits_bits,
  input         io_data_1_in_13_valid,
  input         io_data_1_in_13_bits_valid,
  input  [15:0] io_data_1_in_13_bits_bits,
  input         io_data_1_in_14_valid,
  input         io_data_1_in_14_bits_valid,
  input  [15:0] io_data_1_in_14_bits_bits,
  input         io_data_1_in_15_valid,
  input         io_data_1_in_15_bits_valid,
  input  [15:0] io_data_1_in_15_bits_bits,
  output        io_data_0_out_0_valid,
  output [15:0] io_data_0_out_0_bits,
  output        io_data_0_out_1_valid,
  output [15:0] io_data_0_out_1_bits,
  output        io_data_0_out_2_valid,
  output [15:0] io_data_0_out_2_bits,
  output        io_data_0_out_3_valid,
  output [15:0] io_data_0_out_3_bits,
  output        io_data_0_out_4_valid,
  output [15:0] io_data_0_out_4_bits,
  output        io_data_0_out_5_valid,
  output [15:0] io_data_0_out_5_bits,
  output        io_data_0_out_6_valid,
  output [15:0] io_data_0_out_6_bits,
  output        io_data_0_out_7_valid,
  output [15:0] io_data_0_out_7_bits,
  output        io_data_0_out_8_valid,
  output [15:0] io_data_0_out_8_bits,
  output        io_data_0_out_9_valid,
  output [15:0] io_data_0_out_9_bits,
  output        io_data_0_out_10_valid,
  output [15:0] io_data_0_out_10_bits,
  output        io_data_0_out_11_valid,
  output [15:0] io_data_0_out_11_bits,
  output        io_data_0_out_12_valid,
  output [15:0] io_data_0_out_12_bits,
  output        io_data_0_out_13_valid,
  output [15:0] io_data_0_out_13_bits,
  output        io_data_0_out_14_valid,
  output [15:0] io_data_0_out_14_bits,
  output        io_data_0_out_15_valid,
  output [15:0] io_data_0_out_15_bits,
  input         io_exec_valid,
  input         io_out_valid
);
  wire  MultiDimTime_clock; // @[pearray.scala 63:25]
  wire  MultiDimTime_reset; // @[pearray.scala 63:25]
  wire  MultiDimTime_io_in; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_0; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_1; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_2; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_3; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_4; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_0; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_1; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_2; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_3; // @[pearray.scala 63:25]
  wire  PE_clock; // @[pearray.scala 103:13]
  wire  PE_reset; // @[pearray.scala 103:13]
  wire  PE_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_1_clock; // @[pearray.scala 103:13]
  wire  PE_1_reset; // @[pearray.scala 103:13]
  wire  PE_1_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_2_clock; // @[pearray.scala 103:13]
  wire  PE_2_reset; // @[pearray.scala 103:13]
  wire  PE_2_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_3_clock; // @[pearray.scala 103:13]
  wire  PE_3_reset; // @[pearray.scala 103:13]
  wire  PE_3_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_4_clock; // @[pearray.scala 103:13]
  wire  PE_4_reset; // @[pearray.scala 103:13]
  wire  PE_4_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_5_clock; // @[pearray.scala 103:13]
  wire  PE_5_reset; // @[pearray.scala 103:13]
  wire  PE_5_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_6_clock; // @[pearray.scala 103:13]
  wire  PE_6_reset; // @[pearray.scala 103:13]
  wire  PE_6_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_7_clock; // @[pearray.scala 103:13]
  wire  PE_7_reset; // @[pearray.scala 103:13]
  wire  PE_7_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_8_clock; // @[pearray.scala 103:13]
  wire  PE_8_reset; // @[pearray.scala 103:13]
  wire  PE_8_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_9_clock; // @[pearray.scala 103:13]
  wire  PE_9_reset; // @[pearray.scala 103:13]
  wire  PE_9_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_10_clock; // @[pearray.scala 103:13]
  wire  PE_10_reset; // @[pearray.scala 103:13]
  wire  PE_10_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_11_clock; // @[pearray.scala 103:13]
  wire  PE_11_reset; // @[pearray.scala 103:13]
  wire  PE_11_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_12_clock; // @[pearray.scala 103:13]
  wire  PE_12_reset; // @[pearray.scala 103:13]
  wire  PE_12_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_13_clock; // @[pearray.scala 103:13]
  wire  PE_13_reset; // @[pearray.scala 103:13]
  wire  PE_13_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_14_clock; // @[pearray.scala 103:13]
  wire  PE_14_reset; // @[pearray.scala 103:13]
  wire  PE_14_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_15_clock; // @[pearray.scala 103:13]
  wire  PE_15_reset; // @[pearray.scala 103:13]
  wire  PE_15_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_16_clock; // @[pearray.scala 103:13]
  wire  PE_16_reset; // @[pearray.scala 103:13]
  wire  PE_16_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_17_clock; // @[pearray.scala 103:13]
  wire  PE_17_reset; // @[pearray.scala 103:13]
  wire  PE_17_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_18_clock; // @[pearray.scala 103:13]
  wire  PE_18_reset; // @[pearray.scala 103:13]
  wire  PE_18_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_19_clock; // @[pearray.scala 103:13]
  wire  PE_19_reset; // @[pearray.scala 103:13]
  wire  PE_19_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_20_clock; // @[pearray.scala 103:13]
  wire  PE_20_reset; // @[pearray.scala 103:13]
  wire  PE_20_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_21_clock; // @[pearray.scala 103:13]
  wire  PE_21_reset; // @[pearray.scala 103:13]
  wire  PE_21_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_22_clock; // @[pearray.scala 103:13]
  wire  PE_22_reset; // @[pearray.scala 103:13]
  wire  PE_22_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_23_clock; // @[pearray.scala 103:13]
  wire  PE_23_reset; // @[pearray.scala 103:13]
  wire  PE_23_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_24_clock; // @[pearray.scala 103:13]
  wire  PE_24_reset; // @[pearray.scala 103:13]
  wire  PE_24_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_25_clock; // @[pearray.scala 103:13]
  wire  PE_25_reset; // @[pearray.scala 103:13]
  wire  PE_25_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_26_clock; // @[pearray.scala 103:13]
  wire  PE_26_reset; // @[pearray.scala 103:13]
  wire  PE_26_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_27_clock; // @[pearray.scala 103:13]
  wire  PE_27_reset; // @[pearray.scala 103:13]
  wire  PE_27_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_28_clock; // @[pearray.scala 103:13]
  wire  PE_28_reset; // @[pearray.scala 103:13]
  wire  PE_28_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_29_clock; // @[pearray.scala 103:13]
  wire  PE_29_reset; // @[pearray.scala 103:13]
  wire  PE_29_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_30_clock; // @[pearray.scala 103:13]
  wire  PE_30_reset; // @[pearray.scala 103:13]
  wire  PE_30_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_31_clock; // @[pearray.scala 103:13]
  wire  PE_31_reset; // @[pearray.scala 103:13]
  wire  PE_31_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_32_clock; // @[pearray.scala 103:13]
  wire  PE_32_reset; // @[pearray.scala 103:13]
  wire  PE_32_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_33_clock; // @[pearray.scala 103:13]
  wire  PE_33_reset; // @[pearray.scala 103:13]
  wire  PE_33_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_34_clock; // @[pearray.scala 103:13]
  wire  PE_34_reset; // @[pearray.scala 103:13]
  wire  PE_34_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_35_clock; // @[pearray.scala 103:13]
  wire  PE_35_reset; // @[pearray.scala 103:13]
  wire  PE_35_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_36_clock; // @[pearray.scala 103:13]
  wire  PE_36_reset; // @[pearray.scala 103:13]
  wire  PE_36_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_37_clock; // @[pearray.scala 103:13]
  wire  PE_37_reset; // @[pearray.scala 103:13]
  wire  PE_37_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_38_clock; // @[pearray.scala 103:13]
  wire  PE_38_reset; // @[pearray.scala 103:13]
  wire  PE_38_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_39_clock; // @[pearray.scala 103:13]
  wire  PE_39_reset; // @[pearray.scala 103:13]
  wire  PE_39_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_40_clock; // @[pearray.scala 103:13]
  wire  PE_40_reset; // @[pearray.scala 103:13]
  wire  PE_40_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_41_clock; // @[pearray.scala 103:13]
  wire  PE_41_reset; // @[pearray.scala 103:13]
  wire  PE_41_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_42_clock; // @[pearray.scala 103:13]
  wire  PE_42_reset; // @[pearray.scala 103:13]
  wire  PE_42_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_43_clock; // @[pearray.scala 103:13]
  wire  PE_43_reset; // @[pearray.scala 103:13]
  wire  PE_43_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_44_clock; // @[pearray.scala 103:13]
  wire  PE_44_reset; // @[pearray.scala 103:13]
  wire  PE_44_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_45_clock; // @[pearray.scala 103:13]
  wire  PE_45_reset; // @[pearray.scala 103:13]
  wire  PE_45_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_46_clock; // @[pearray.scala 103:13]
  wire  PE_46_reset; // @[pearray.scala 103:13]
  wire  PE_46_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_47_clock; // @[pearray.scala 103:13]
  wire  PE_47_reset; // @[pearray.scala 103:13]
  wire  PE_47_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_48_clock; // @[pearray.scala 103:13]
  wire  PE_48_reset; // @[pearray.scala 103:13]
  wire  PE_48_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_49_clock; // @[pearray.scala 103:13]
  wire  PE_49_reset; // @[pearray.scala 103:13]
  wire  PE_49_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_50_clock; // @[pearray.scala 103:13]
  wire  PE_50_reset; // @[pearray.scala 103:13]
  wire  PE_50_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_51_clock; // @[pearray.scala 103:13]
  wire  PE_51_reset; // @[pearray.scala 103:13]
  wire  PE_51_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_52_clock; // @[pearray.scala 103:13]
  wire  PE_52_reset; // @[pearray.scala 103:13]
  wire  PE_52_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_53_clock; // @[pearray.scala 103:13]
  wire  PE_53_reset; // @[pearray.scala 103:13]
  wire  PE_53_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_54_clock; // @[pearray.scala 103:13]
  wire  PE_54_reset; // @[pearray.scala 103:13]
  wire  PE_54_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_55_clock; // @[pearray.scala 103:13]
  wire  PE_55_reset; // @[pearray.scala 103:13]
  wire  PE_55_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_56_clock; // @[pearray.scala 103:13]
  wire  PE_56_reset; // @[pearray.scala 103:13]
  wire  PE_56_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_57_clock; // @[pearray.scala 103:13]
  wire  PE_57_reset; // @[pearray.scala 103:13]
  wire  PE_57_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_58_clock; // @[pearray.scala 103:13]
  wire  PE_58_reset; // @[pearray.scala 103:13]
  wire  PE_58_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_59_clock; // @[pearray.scala 103:13]
  wire  PE_59_reset; // @[pearray.scala 103:13]
  wire  PE_59_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_60_clock; // @[pearray.scala 103:13]
  wire  PE_60_reset; // @[pearray.scala 103:13]
  wire  PE_60_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_61_clock; // @[pearray.scala 103:13]
  wire  PE_61_reset; // @[pearray.scala 103:13]
  wire  PE_61_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_62_clock; // @[pearray.scala 103:13]
  wire  PE_62_reset; // @[pearray.scala 103:13]
  wire  PE_62_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_63_clock; // @[pearray.scala 103:13]
  wire  PE_63_reset; // @[pearray.scala 103:13]
  wire  PE_63_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_64_clock; // @[pearray.scala 103:13]
  wire  PE_64_reset; // @[pearray.scala 103:13]
  wire  PE_64_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_64_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_64_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_64_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_64_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_64_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_64_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_64_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_64_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_64_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_64_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_64_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_64_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_65_clock; // @[pearray.scala 103:13]
  wire  PE_65_reset; // @[pearray.scala 103:13]
  wire  PE_65_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_65_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_65_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_65_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_65_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_65_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_65_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_65_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_65_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_65_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_65_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_65_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_65_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_66_clock; // @[pearray.scala 103:13]
  wire  PE_66_reset; // @[pearray.scala 103:13]
  wire  PE_66_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_66_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_66_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_66_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_66_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_66_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_66_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_66_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_66_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_66_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_66_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_66_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_66_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_67_clock; // @[pearray.scala 103:13]
  wire  PE_67_reset; // @[pearray.scala 103:13]
  wire  PE_67_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_67_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_67_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_67_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_67_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_67_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_67_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_67_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_67_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_67_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_67_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_67_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_67_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_68_clock; // @[pearray.scala 103:13]
  wire  PE_68_reset; // @[pearray.scala 103:13]
  wire  PE_68_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_68_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_68_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_68_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_68_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_68_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_68_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_68_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_68_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_68_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_68_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_68_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_68_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_69_clock; // @[pearray.scala 103:13]
  wire  PE_69_reset; // @[pearray.scala 103:13]
  wire  PE_69_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_69_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_69_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_69_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_69_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_69_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_69_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_69_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_69_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_69_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_69_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_69_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_69_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_70_clock; // @[pearray.scala 103:13]
  wire  PE_70_reset; // @[pearray.scala 103:13]
  wire  PE_70_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_70_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_70_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_70_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_70_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_70_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_70_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_70_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_70_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_70_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_70_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_70_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_70_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_71_clock; // @[pearray.scala 103:13]
  wire  PE_71_reset; // @[pearray.scala 103:13]
  wire  PE_71_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_71_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_71_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_71_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_71_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_71_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_71_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_71_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_71_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_71_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_71_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_71_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_71_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_72_clock; // @[pearray.scala 103:13]
  wire  PE_72_reset; // @[pearray.scala 103:13]
  wire  PE_72_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_72_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_72_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_72_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_72_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_72_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_72_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_72_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_72_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_72_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_72_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_72_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_72_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_73_clock; // @[pearray.scala 103:13]
  wire  PE_73_reset; // @[pearray.scala 103:13]
  wire  PE_73_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_73_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_73_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_73_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_73_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_73_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_73_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_73_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_73_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_73_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_73_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_73_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_73_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_74_clock; // @[pearray.scala 103:13]
  wire  PE_74_reset; // @[pearray.scala 103:13]
  wire  PE_74_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_74_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_74_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_74_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_74_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_74_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_74_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_74_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_74_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_74_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_74_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_74_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_74_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_75_clock; // @[pearray.scala 103:13]
  wire  PE_75_reset; // @[pearray.scala 103:13]
  wire  PE_75_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_75_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_75_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_75_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_75_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_75_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_75_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_75_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_75_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_75_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_75_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_75_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_75_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_76_clock; // @[pearray.scala 103:13]
  wire  PE_76_reset; // @[pearray.scala 103:13]
  wire  PE_76_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_76_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_76_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_76_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_76_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_76_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_76_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_76_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_76_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_76_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_76_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_76_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_76_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_77_clock; // @[pearray.scala 103:13]
  wire  PE_77_reset; // @[pearray.scala 103:13]
  wire  PE_77_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_77_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_77_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_77_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_77_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_77_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_77_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_77_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_77_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_77_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_77_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_77_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_77_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_78_clock; // @[pearray.scala 103:13]
  wire  PE_78_reset; // @[pearray.scala 103:13]
  wire  PE_78_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_78_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_78_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_78_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_78_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_78_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_78_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_78_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_78_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_78_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_78_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_78_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_78_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_79_clock; // @[pearray.scala 103:13]
  wire  PE_79_reset; // @[pearray.scala 103:13]
  wire  PE_79_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_79_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_79_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_79_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_79_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_79_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_79_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_79_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_79_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_79_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_79_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_79_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_79_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_80_clock; // @[pearray.scala 103:13]
  wire  PE_80_reset; // @[pearray.scala 103:13]
  wire  PE_80_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_80_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_80_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_80_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_80_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_80_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_80_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_80_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_80_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_80_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_80_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_80_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_80_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_81_clock; // @[pearray.scala 103:13]
  wire  PE_81_reset; // @[pearray.scala 103:13]
  wire  PE_81_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_81_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_81_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_81_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_81_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_81_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_81_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_81_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_81_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_81_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_81_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_81_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_81_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_82_clock; // @[pearray.scala 103:13]
  wire  PE_82_reset; // @[pearray.scala 103:13]
  wire  PE_82_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_82_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_82_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_82_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_82_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_82_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_82_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_82_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_82_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_82_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_82_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_82_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_82_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_83_clock; // @[pearray.scala 103:13]
  wire  PE_83_reset; // @[pearray.scala 103:13]
  wire  PE_83_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_83_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_83_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_83_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_83_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_83_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_83_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_83_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_83_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_83_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_83_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_83_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_83_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_84_clock; // @[pearray.scala 103:13]
  wire  PE_84_reset; // @[pearray.scala 103:13]
  wire  PE_84_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_84_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_84_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_84_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_84_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_84_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_84_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_84_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_84_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_84_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_84_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_84_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_84_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_85_clock; // @[pearray.scala 103:13]
  wire  PE_85_reset; // @[pearray.scala 103:13]
  wire  PE_85_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_85_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_85_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_85_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_85_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_85_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_85_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_85_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_85_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_85_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_85_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_85_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_85_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_86_clock; // @[pearray.scala 103:13]
  wire  PE_86_reset; // @[pearray.scala 103:13]
  wire  PE_86_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_86_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_86_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_86_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_86_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_86_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_86_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_86_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_86_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_86_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_86_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_86_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_86_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_87_clock; // @[pearray.scala 103:13]
  wire  PE_87_reset; // @[pearray.scala 103:13]
  wire  PE_87_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_87_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_87_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_87_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_87_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_87_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_87_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_87_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_87_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_87_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_87_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_87_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_87_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_88_clock; // @[pearray.scala 103:13]
  wire  PE_88_reset; // @[pearray.scala 103:13]
  wire  PE_88_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_88_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_88_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_88_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_88_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_88_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_88_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_88_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_88_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_88_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_88_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_88_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_88_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_89_clock; // @[pearray.scala 103:13]
  wire  PE_89_reset; // @[pearray.scala 103:13]
  wire  PE_89_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_89_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_89_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_89_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_89_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_89_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_89_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_89_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_89_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_89_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_89_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_89_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_89_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_90_clock; // @[pearray.scala 103:13]
  wire  PE_90_reset; // @[pearray.scala 103:13]
  wire  PE_90_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_90_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_90_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_90_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_90_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_90_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_90_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_90_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_90_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_90_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_90_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_90_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_90_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_91_clock; // @[pearray.scala 103:13]
  wire  PE_91_reset; // @[pearray.scala 103:13]
  wire  PE_91_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_91_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_91_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_91_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_91_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_91_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_91_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_91_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_91_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_91_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_91_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_91_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_91_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_92_clock; // @[pearray.scala 103:13]
  wire  PE_92_reset; // @[pearray.scala 103:13]
  wire  PE_92_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_92_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_92_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_92_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_92_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_92_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_92_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_92_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_92_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_92_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_92_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_92_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_92_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_93_clock; // @[pearray.scala 103:13]
  wire  PE_93_reset; // @[pearray.scala 103:13]
  wire  PE_93_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_93_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_93_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_93_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_93_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_93_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_93_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_93_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_93_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_93_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_93_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_93_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_93_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_94_clock; // @[pearray.scala 103:13]
  wire  PE_94_reset; // @[pearray.scala 103:13]
  wire  PE_94_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_94_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_94_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_94_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_94_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_94_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_94_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_94_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_94_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_94_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_94_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_94_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_94_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_95_clock; // @[pearray.scala 103:13]
  wire  PE_95_reset; // @[pearray.scala 103:13]
  wire  PE_95_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_95_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_95_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_95_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_95_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_95_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_95_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_95_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_95_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_95_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_95_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_95_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_95_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_96_clock; // @[pearray.scala 103:13]
  wire  PE_96_reset; // @[pearray.scala 103:13]
  wire  PE_96_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_96_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_96_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_96_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_96_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_96_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_96_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_96_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_96_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_96_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_96_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_96_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_96_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_97_clock; // @[pearray.scala 103:13]
  wire  PE_97_reset; // @[pearray.scala 103:13]
  wire  PE_97_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_97_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_97_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_97_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_97_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_97_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_97_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_97_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_97_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_97_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_97_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_97_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_97_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_98_clock; // @[pearray.scala 103:13]
  wire  PE_98_reset; // @[pearray.scala 103:13]
  wire  PE_98_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_98_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_98_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_98_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_98_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_98_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_98_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_98_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_98_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_98_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_98_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_98_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_98_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_99_clock; // @[pearray.scala 103:13]
  wire  PE_99_reset; // @[pearray.scala 103:13]
  wire  PE_99_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_99_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_99_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_99_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_99_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_99_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_99_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_99_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_99_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_99_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_99_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_99_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_99_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_100_clock; // @[pearray.scala 103:13]
  wire  PE_100_reset; // @[pearray.scala 103:13]
  wire  PE_100_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_100_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_100_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_100_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_100_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_100_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_100_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_100_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_100_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_100_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_100_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_100_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_100_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_101_clock; // @[pearray.scala 103:13]
  wire  PE_101_reset; // @[pearray.scala 103:13]
  wire  PE_101_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_101_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_101_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_101_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_101_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_101_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_101_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_101_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_101_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_101_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_101_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_101_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_101_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_102_clock; // @[pearray.scala 103:13]
  wire  PE_102_reset; // @[pearray.scala 103:13]
  wire  PE_102_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_102_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_102_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_102_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_102_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_102_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_102_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_102_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_102_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_102_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_102_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_102_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_102_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_103_clock; // @[pearray.scala 103:13]
  wire  PE_103_reset; // @[pearray.scala 103:13]
  wire  PE_103_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_103_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_103_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_103_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_103_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_103_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_103_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_103_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_103_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_103_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_103_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_103_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_103_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_104_clock; // @[pearray.scala 103:13]
  wire  PE_104_reset; // @[pearray.scala 103:13]
  wire  PE_104_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_104_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_104_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_104_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_104_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_104_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_104_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_104_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_104_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_104_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_104_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_104_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_104_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_105_clock; // @[pearray.scala 103:13]
  wire  PE_105_reset; // @[pearray.scala 103:13]
  wire  PE_105_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_105_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_105_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_105_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_105_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_105_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_105_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_105_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_105_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_105_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_105_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_105_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_105_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_106_clock; // @[pearray.scala 103:13]
  wire  PE_106_reset; // @[pearray.scala 103:13]
  wire  PE_106_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_106_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_106_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_106_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_106_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_106_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_106_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_106_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_106_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_106_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_106_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_106_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_106_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_107_clock; // @[pearray.scala 103:13]
  wire  PE_107_reset; // @[pearray.scala 103:13]
  wire  PE_107_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_107_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_107_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_107_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_107_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_107_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_107_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_107_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_107_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_107_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_107_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_107_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_107_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_108_clock; // @[pearray.scala 103:13]
  wire  PE_108_reset; // @[pearray.scala 103:13]
  wire  PE_108_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_108_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_108_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_108_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_108_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_108_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_108_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_108_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_108_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_108_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_108_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_108_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_108_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_109_clock; // @[pearray.scala 103:13]
  wire  PE_109_reset; // @[pearray.scala 103:13]
  wire  PE_109_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_109_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_109_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_109_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_109_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_109_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_109_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_109_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_109_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_109_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_109_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_109_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_109_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_110_clock; // @[pearray.scala 103:13]
  wire  PE_110_reset; // @[pearray.scala 103:13]
  wire  PE_110_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_110_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_110_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_110_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_110_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_110_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_110_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_110_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_110_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_110_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_110_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_110_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_110_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_111_clock; // @[pearray.scala 103:13]
  wire  PE_111_reset; // @[pearray.scala 103:13]
  wire  PE_111_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_111_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_111_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_111_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_111_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_111_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_111_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_111_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_111_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_111_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_111_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_111_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_111_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_112_clock; // @[pearray.scala 103:13]
  wire  PE_112_reset; // @[pearray.scala 103:13]
  wire  PE_112_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_112_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_112_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_112_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_112_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_112_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_112_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_112_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_112_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_112_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_112_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_112_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_112_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_113_clock; // @[pearray.scala 103:13]
  wire  PE_113_reset; // @[pearray.scala 103:13]
  wire  PE_113_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_113_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_113_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_113_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_113_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_113_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_113_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_113_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_113_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_113_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_113_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_113_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_113_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_114_clock; // @[pearray.scala 103:13]
  wire  PE_114_reset; // @[pearray.scala 103:13]
  wire  PE_114_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_114_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_114_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_114_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_114_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_114_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_114_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_114_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_114_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_114_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_114_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_114_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_114_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_115_clock; // @[pearray.scala 103:13]
  wire  PE_115_reset; // @[pearray.scala 103:13]
  wire  PE_115_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_115_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_115_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_115_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_115_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_115_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_115_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_115_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_115_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_115_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_115_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_115_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_115_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_116_clock; // @[pearray.scala 103:13]
  wire  PE_116_reset; // @[pearray.scala 103:13]
  wire  PE_116_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_116_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_116_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_116_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_116_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_116_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_116_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_116_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_116_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_116_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_116_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_116_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_116_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_117_clock; // @[pearray.scala 103:13]
  wire  PE_117_reset; // @[pearray.scala 103:13]
  wire  PE_117_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_117_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_117_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_117_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_117_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_117_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_117_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_117_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_117_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_117_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_117_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_117_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_117_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_118_clock; // @[pearray.scala 103:13]
  wire  PE_118_reset; // @[pearray.scala 103:13]
  wire  PE_118_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_118_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_118_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_118_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_118_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_118_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_118_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_118_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_118_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_118_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_118_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_118_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_118_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_119_clock; // @[pearray.scala 103:13]
  wire  PE_119_reset; // @[pearray.scala 103:13]
  wire  PE_119_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_119_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_119_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_119_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_119_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_119_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_119_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_119_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_119_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_119_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_119_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_119_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_119_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_120_clock; // @[pearray.scala 103:13]
  wire  PE_120_reset; // @[pearray.scala 103:13]
  wire  PE_120_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_120_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_120_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_120_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_120_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_120_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_120_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_120_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_120_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_120_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_120_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_120_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_120_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_121_clock; // @[pearray.scala 103:13]
  wire  PE_121_reset; // @[pearray.scala 103:13]
  wire  PE_121_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_121_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_121_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_121_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_121_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_121_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_121_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_121_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_121_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_121_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_121_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_121_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_121_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_122_clock; // @[pearray.scala 103:13]
  wire  PE_122_reset; // @[pearray.scala 103:13]
  wire  PE_122_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_122_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_122_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_122_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_122_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_122_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_122_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_122_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_122_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_122_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_122_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_122_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_122_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_123_clock; // @[pearray.scala 103:13]
  wire  PE_123_reset; // @[pearray.scala 103:13]
  wire  PE_123_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_123_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_123_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_123_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_123_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_123_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_123_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_123_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_123_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_123_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_123_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_123_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_123_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_124_clock; // @[pearray.scala 103:13]
  wire  PE_124_reset; // @[pearray.scala 103:13]
  wire  PE_124_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_124_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_124_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_124_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_124_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_124_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_124_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_124_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_124_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_124_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_124_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_124_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_124_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_125_clock; // @[pearray.scala 103:13]
  wire  PE_125_reset; // @[pearray.scala 103:13]
  wire  PE_125_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_125_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_125_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_125_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_125_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_125_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_125_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_125_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_125_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_125_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_125_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_125_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_125_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_126_clock; // @[pearray.scala 103:13]
  wire  PE_126_reset; // @[pearray.scala 103:13]
  wire  PE_126_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_126_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_126_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_126_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_126_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_126_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_126_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_126_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_126_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_126_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_126_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_126_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_126_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_127_clock; // @[pearray.scala 103:13]
  wire  PE_127_reset; // @[pearray.scala 103:13]
  wire  PE_127_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_127_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_127_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_127_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_127_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_127_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_127_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_127_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_127_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_127_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_127_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_127_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_127_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_128_clock; // @[pearray.scala 103:13]
  wire  PE_128_reset; // @[pearray.scala 103:13]
  wire  PE_128_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_128_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_128_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_128_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_128_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_128_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_128_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_128_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_128_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_128_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_128_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_128_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_128_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_129_clock; // @[pearray.scala 103:13]
  wire  PE_129_reset; // @[pearray.scala 103:13]
  wire  PE_129_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_129_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_129_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_129_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_129_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_129_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_129_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_129_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_129_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_129_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_129_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_129_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_129_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_130_clock; // @[pearray.scala 103:13]
  wire  PE_130_reset; // @[pearray.scala 103:13]
  wire  PE_130_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_130_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_130_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_130_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_130_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_130_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_130_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_130_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_130_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_130_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_130_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_130_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_130_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_131_clock; // @[pearray.scala 103:13]
  wire  PE_131_reset; // @[pearray.scala 103:13]
  wire  PE_131_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_131_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_131_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_131_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_131_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_131_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_131_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_131_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_131_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_131_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_131_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_131_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_131_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_132_clock; // @[pearray.scala 103:13]
  wire  PE_132_reset; // @[pearray.scala 103:13]
  wire  PE_132_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_132_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_132_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_132_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_132_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_132_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_132_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_132_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_132_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_132_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_132_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_132_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_132_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_133_clock; // @[pearray.scala 103:13]
  wire  PE_133_reset; // @[pearray.scala 103:13]
  wire  PE_133_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_133_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_133_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_133_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_133_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_133_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_133_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_133_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_133_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_133_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_133_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_133_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_133_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_134_clock; // @[pearray.scala 103:13]
  wire  PE_134_reset; // @[pearray.scala 103:13]
  wire  PE_134_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_134_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_134_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_134_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_134_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_134_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_134_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_134_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_134_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_134_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_134_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_134_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_134_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_135_clock; // @[pearray.scala 103:13]
  wire  PE_135_reset; // @[pearray.scala 103:13]
  wire  PE_135_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_135_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_135_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_135_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_135_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_135_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_135_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_135_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_135_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_135_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_135_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_135_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_135_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_136_clock; // @[pearray.scala 103:13]
  wire  PE_136_reset; // @[pearray.scala 103:13]
  wire  PE_136_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_136_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_136_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_136_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_136_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_136_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_136_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_136_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_136_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_136_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_136_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_136_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_136_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_137_clock; // @[pearray.scala 103:13]
  wire  PE_137_reset; // @[pearray.scala 103:13]
  wire  PE_137_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_137_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_137_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_137_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_137_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_137_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_137_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_137_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_137_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_137_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_137_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_137_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_137_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_138_clock; // @[pearray.scala 103:13]
  wire  PE_138_reset; // @[pearray.scala 103:13]
  wire  PE_138_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_138_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_138_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_138_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_138_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_138_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_138_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_138_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_138_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_138_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_138_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_138_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_138_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_139_clock; // @[pearray.scala 103:13]
  wire  PE_139_reset; // @[pearray.scala 103:13]
  wire  PE_139_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_139_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_139_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_139_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_139_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_139_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_139_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_139_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_139_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_139_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_139_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_139_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_139_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_140_clock; // @[pearray.scala 103:13]
  wire  PE_140_reset; // @[pearray.scala 103:13]
  wire  PE_140_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_140_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_140_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_140_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_140_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_140_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_140_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_140_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_140_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_140_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_140_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_140_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_140_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_141_clock; // @[pearray.scala 103:13]
  wire  PE_141_reset; // @[pearray.scala 103:13]
  wire  PE_141_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_141_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_141_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_141_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_141_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_141_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_141_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_141_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_141_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_141_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_141_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_141_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_141_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_142_clock; // @[pearray.scala 103:13]
  wire  PE_142_reset; // @[pearray.scala 103:13]
  wire  PE_142_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_142_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_142_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_142_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_142_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_142_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_142_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_142_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_142_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_142_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_142_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_142_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_142_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_143_clock; // @[pearray.scala 103:13]
  wire  PE_143_reset; // @[pearray.scala 103:13]
  wire  PE_143_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_143_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_143_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_143_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_143_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_143_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_143_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_143_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_143_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_143_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_143_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_143_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_143_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_144_clock; // @[pearray.scala 103:13]
  wire  PE_144_reset; // @[pearray.scala 103:13]
  wire  PE_144_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_144_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_144_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_144_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_144_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_144_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_144_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_144_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_144_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_144_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_144_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_144_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_144_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_145_clock; // @[pearray.scala 103:13]
  wire  PE_145_reset; // @[pearray.scala 103:13]
  wire  PE_145_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_145_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_145_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_145_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_145_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_145_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_145_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_145_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_145_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_145_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_145_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_145_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_145_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_146_clock; // @[pearray.scala 103:13]
  wire  PE_146_reset; // @[pearray.scala 103:13]
  wire  PE_146_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_146_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_146_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_146_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_146_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_146_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_146_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_146_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_146_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_146_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_146_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_146_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_146_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_147_clock; // @[pearray.scala 103:13]
  wire  PE_147_reset; // @[pearray.scala 103:13]
  wire  PE_147_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_147_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_147_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_147_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_147_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_147_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_147_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_147_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_147_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_147_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_147_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_147_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_147_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_148_clock; // @[pearray.scala 103:13]
  wire  PE_148_reset; // @[pearray.scala 103:13]
  wire  PE_148_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_148_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_148_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_148_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_148_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_148_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_148_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_148_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_148_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_148_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_148_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_148_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_148_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_149_clock; // @[pearray.scala 103:13]
  wire  PE_149_reset; // @[pearray.scala 103:13]
  wire  PE_149_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_149_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_149_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_149_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_149_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_149_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_149_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_149_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_149_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_149_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_149_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_149_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_149_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_150_clock; // @[pearray.scala 103:13]
  wire  PE_150_reset; // @[pearray.scala 103:13]
  wire  PE_150_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_150_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_150_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_150_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_150_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_150_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_150_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_150_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_150_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_150_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_150_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_150_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_150_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_151_clock; // @[pearray.scala 103:13]
  wire  PE_151_reset; // @[pearray.scala 103:13]
  wire  PE_151_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_151_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_151_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_151_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_151_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_151_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_151_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_151_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_151_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_151_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_151_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_151_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_151_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_152_clock; // @[pearray.scala 103:13]
  wire  PE_152_reset; // @[pearray.scala 103:13]
  wire  PE_152_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_152_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_152_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_152_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_152_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_152_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_152_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_152_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_152_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_152_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_152_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_152_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_152_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_153_clock; // @[pearray.scala 103:13]
  wire  PE_153_reset; // @[pearray.scala 103:13]
  wire  PE_153_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_153_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_153_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_153_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_153_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_153_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_153_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_153_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_153_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_153_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_153_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_153_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_153_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_154_clock; // @[pearray.scala 103:13]
  wire  PE_154_reset; // @[pearray.scala 103:13]
  wire  PE_154_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_154_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_154_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_154_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_154_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_154_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_154_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_154_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_154_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_154_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_154_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_154_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_154_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_155_clock; // @[pearray.scala 103:13]
  wire  PE_155_reset; // @[pearray.scala 103:13]
  wire  PE_155_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_155_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_155_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_155_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_155_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_155_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_155_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_155_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_155_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_155_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_155_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_155_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_155_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_156_clock; // @[pearray.scala 103:13]
  wire  PE_156_reset; // @[pearray.scala 103:13]
  wire  PE_156_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_156_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_156_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_156_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_156_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_156_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_156_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_156_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_156_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_156_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_156_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_156_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_156_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_157_clock; // @[pearray.scala 103:13]
  wire  PE_157_reset; // @[pearray.scala 103:13]
  wire  PE_157_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_157_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_157_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_157_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_157_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_157_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_157_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_157_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_157_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_157_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_157_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_157_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_157_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_158_clock; // @[pearray.scala 103:13]
  wire  PE_158_reset; // @[pearray.scala 103:13]
  wire  PE_158_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_158_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_158_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_158_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_158_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_158_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_158_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_158_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_158_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_158_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_158_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_158_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_158_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_159_clock; // @[pearray.scala 103:13]
  wire  PE_159_reset; // @[pearray.scala 103:13]
  wire  PE_159_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_159_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_159_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_159_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_159_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_159_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_159_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_159_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_159_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_159_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_159_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_159_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_159_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_160_clock; // @[pearray.scala 103:13]
  wire  PE_160_reset; // @[pearray.scala 103:13]
  wire  PE_160_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_160_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_160_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_160_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_160_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_160_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_160_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_160_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_160_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_160_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_160_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_160_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_160_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_161_clock; // @[pearray.scala 103:13]
  wire  PE_161_reset; // @[pearray.scala 103:13]
  wire  PE_161_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_161_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_161_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_161_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_161_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_161_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_161_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_161_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_161_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_161_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_161_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_161_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_161_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_162_clock; // @[pearray.scala 103:13]
  wire  PE_162_reset; // @[pearray.scala 103:13]
  wire  PE_162_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_162_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_162_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_162_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_162_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_162_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_162_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_162_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_162_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_162_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_162_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_162_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_162_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_163_clock; // @[pearray.scala 103:13]
  wire  PE_163_reset; // @[pearray.scala 103:13]
  wire  PE_163_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_163_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_163_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_163_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_163_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_163_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_163_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_163_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_163_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_163_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_163_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_163_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_163_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_164_clock; // @[pearray.scala 103:13]
  wire  PE_164_reset; // @[pearray.scala 103:13]
  wire  PE_164_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_164_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_164_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_164_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_164_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_164_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_164_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_164_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_164_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_164_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_164_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_164_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_164_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_165_clock; // @[pearray.scala 103:13]
  wire  PE_165_reset; // @[pearray.scala 103:13]
  wire  PE_165_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_165_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_165_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_165_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_165_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_165_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_165_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_165_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_165_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_165_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_165_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_165_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_165_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_166_clock; // @[pearray.scala 103:13]
  wire  PE_166_reset; // @[pearray.scala 103:13]
  wire  PE_166_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_166_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_166_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_166_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_166_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_166_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_166_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_166_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_166_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_166_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_166_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_166_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_166_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_167_clock; // @[pearray.scala 103:13]
  wire  PE_167_reset; // @[pearray.scala 103:13]
  wire  PE_167_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_167_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_167_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_167_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_167_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_167_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_167_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_167_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_167_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_167_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_167_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_167_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_167_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_168_clock; // @[pearray.scala 103:13]
  wire  PE_168_reset; // @[pearray.scala 103:13]
  wire  PE_168_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_168_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_168_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_168_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_168_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_168_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_168_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_168_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_168_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_168_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_168_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_168_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_168_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_169_clock; // @[pearray.scala 103:13]
  wire  PE_169_reset; // @[pearray.scala 103:13]
  wire  PE_169_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_169_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_169_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_169_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_169_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_169_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_169_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_169_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_169_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_169_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_169_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_169_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_169_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_170_clock; // @[pearray.scala 103:13]
  wire  PE_170_reset; // @[pearray.scala 103:13]
  wire  PE_170_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_170_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_170_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_170_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_170_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_170_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_170_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_170_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_170_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_170_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_170_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_170_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_170_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_171_clock; // @[pearray.scala 103:13]
  wire  PE_171_reset; // @[pearray.scala 103:13]
  wire  PE_171_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_171_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_171_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_171_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_171_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_171_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_171_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_171_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_171_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_171_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_171_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_171_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_171_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_172_clock; // @[pearray.scala 103:13]
  wire  PE_172_reset; // @[pearray.scala 103:13]
  wire  PE_172_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_172_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_172_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_172_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_172_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_172_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_172_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_172_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_172_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_172_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_172_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_172_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_172_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_173_clock; // @[pearray.scala 103:13]
  wire  PE_173_reset; // @[pearray.scala 103:13]
  wire  PE_173_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_173_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_173_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_173_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_173_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_173_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_173_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_173_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_173_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_173_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_173_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_173_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_173_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_174_clock; // @[pearray.scala 103:13]
  wire  PE_174_reset; // @[pearray.scala 103:13]
  wire  PE_174_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_174_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_174_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_174_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_174_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_174_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_174_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_174_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_174_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_174_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_174_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_174_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_174_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_175_clock; // @[pearray.scala 103:13]
  wire  PE_175_reset; // @[pearray.scala 103:13]
  wire  PE_175_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_175_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_175_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_175_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_175_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_175_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_175_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_175_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_175_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_175_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_175_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_175_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_175_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_176_clock; // @[pearray.scala 103:13]
  wire  PE_176_reset; // @[pearray.scala 103:13]
  wire  PE_176_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_176_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_176_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_176_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_176_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_176_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_176_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_176_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_176_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_176_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_176_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_176_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_176_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_177_clock; // @[pearray.scala 103:13]
  wire  PE_177_reset; // @[pearray.scala 103:13]
  wire  PE_177_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_177_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_177_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_177_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_177_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_177_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_177_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_177_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_177_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_177_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_177_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_177_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_177_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_178_clock; // @[pearray.scala 103:13]
  wire  PE_178_reset; // @[pearray.scala 103:13]
  wire  PE_178_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_178_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_178_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_178_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_178_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_178_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_178_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_178_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_178_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_178_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_178_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_178_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_178_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_179_clock; // @[pearray.scala 103:13]
  wire  PE_179_reset; // @[pearray.scala 103:13]
  wire  PE_179_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_179_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_179_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_179_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_179_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_179_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_179_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_179_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_179_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_179_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_179_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_179_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_179_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_180_clock; // @[pearray.scala 103:13]
  wire  PE_180_reset; // @[pearray.scala 103:13]
  wire  PE_180_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_180_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_180_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_180_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_180_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_180_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_180_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_180_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_180_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_180_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_180_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_180_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_180_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_181_clock; // @[pearray.scala 103:13]
  wire  PE_181_reset; // @[pearray.scala 103:13]
  wire  PE_181_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_181_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_181_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_181_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_181_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_181_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_181_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_181_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_181_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_181_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_181_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_181_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_181_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_182_clock; // @[pearray.scala 103:13]
  wire  PE_182_reset; // @[pearray.scala 103:13]
  wire  PE_182_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_182_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_182_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_182_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_182_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_182_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_182_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_182_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_182_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_182_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_182_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_182_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_182_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_183_clock; // @[pearray.scala 103:13]
  wire  PE_183_reset; // @[pearray.scala 103:13]
  wire  PE_183_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_183_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_183_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_183_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_183_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_183_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_183_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_183_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_183_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_183_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_183_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_183_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_183_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_184_clock; // @[pearray.scala 103:13]
  wire  PE_184_reset; // @[pearray.scala 103:13]
  wire  PE_184_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_184_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_184_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_184_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_184_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_184_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_184_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_184_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_184_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_184_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_184_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_184_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_184_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_185_clock; // @[pearray.scala 103:13]
  wire  PE_185_reset; // @[pearray.scala 103:13]
  wire  PE_185_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_185_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_185_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_185_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_185_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_185_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_185_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_185_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_185_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_185_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_185_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_185_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_185_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_186_clock; // @[pearray.scala 103:13]
  wire  PE_186_reset; // @[pearray.scala 103:13]
  wire  PE_186_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_186_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_186_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_186_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_186_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_186_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_186_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_186_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_186_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_186_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_186_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_186_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_186_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_187_clock; // @[pearray.scala 103:13]
  wire  PE_187_reset; // @[pearray.scala 103:13]
  wire  PE_187_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_187_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_187_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_187_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_187_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_187_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_187_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_187_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_187_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_187_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_187_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_187_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_187_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_188_clock; // @[pearray.scala 103:13]
  wire  PE_188_reset; // @[pearray.scala 103:13]
  wire  PE_188_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_188_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_188_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_188_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_188_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_188_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_188_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_188_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_188_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_188_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_188_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_188_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_188_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_189_clock; // @[pearray.scala 103:13]
  wire  PE_189_reset; // @[pearray.scala 103:13]
  wire  PE_189_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_189_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_189_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_189_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_189_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_189_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_189_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_189_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_189_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_189_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_189_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_189_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_189_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_190_clock; // @[pearray.scala 103:13]
  wire  PE_190_reset; // @[pearray.scala 103:13]
  wire  PE_190_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_190_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_190_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_190_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_190_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_190_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_190_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_190_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_190_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_190_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_190_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_190_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_190_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_191_clock; // @[pearray.scala 103:13]
  wire  PE_191_reset; // @[pearray.scala 103:13]
  wire  PE_191_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_191_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_191_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_191_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_191_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_191_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_191_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_191_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_191_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_191_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_191_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_191_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_191_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_192_clock; // @[pearray.scala 103:13]
  wire  PE_192_reset; // @[pearray.scala 103:13]
  wire  PE_192_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_192_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_192_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_192_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_192_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_192_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_192_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_192_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_192_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_192_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_192_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_192_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_192_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_193_clock; // @[pearray.scala 103:13]
  wire  PE_193_reset; // @[pearray.scala 103:13]
  wire  PE_193_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_193_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_193_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_193_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_193_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_193_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_193_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_193_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_193_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_193_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_193_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_193_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_193_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_194_clock; // @[pearray.scala 103:13]
  wire  PE_194_reset; // @[pearray.scala 103:13]
  wire  PE_194_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_194_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_194_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_194_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_194_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_194_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_194_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_194_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_194_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_194_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_194_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_194_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_194_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_195_clock; // @[pearray.scala 103:13]
  wire  PE_195_reset; // @[pearray.scala 103:13]
  wire  PE_195_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_195_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_195_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_195_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_195_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_195_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_195_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_195_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_195_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_195_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_195_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_195_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_195_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_196_clock; // @[pearray.scala 103:13]
  wire  PE_196_reset; // @[pearray.scala 103:13]
  wire  PE_196_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_196_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_196_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_196_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_196_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_196_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_196_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_196_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_196_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_196_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_196_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_196_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_196_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_197_clock; // @[pearray.scala 103:13]
  wire  PE_197_reset; // @[pearray.scala 103:13]
  wire  PE_197_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_197_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_197_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_197_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_197_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_197_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_197_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_197_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_197_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_197_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_197_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_197_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_197_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_198_clock; // @[pearray.scala 103:13]
  wire  PE_198_reset; // @[pearray.scala 103:13]
  wire  PE_198_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_198_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_198_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_198_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_198_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_198_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_198_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_198_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_198_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_198_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_198_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_198_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_198_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_199_clock; // @[pearray.scala 103:13]
  wire  PE_199_reset; // @[pearray.scala 103:13]
  wire  PE_199_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_199_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_199_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_199_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_199_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_199_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_199_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_199_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_199_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_199_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_199_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_199_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_199_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_200_clock; // @[pearray.scala 103:13]
  wire  PE_200_reset; // @[pearray.scala 103:13]
  wire  PE_200_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_200_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_200_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_200_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_200_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_200_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_200_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_200_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_200_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_200_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_200_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_200_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_200_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_201_clock; // @[pearray.scala 103:13]
  wire  PE_201_reset; // @[pearray.scala 103:13]
  wire  PE_201_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_201_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_201_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_201_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_201_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_201_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_201_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_201_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_201_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_201_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_201_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_201_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_201_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_202_clock; // @[pearray.scala 103:13]
  wire  PE_202_reset; // @[pearray.scala 103:13]
  wire  PE_202_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_202_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_202_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_202_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_202_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_202_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_202_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_202_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_202_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_202_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_202_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_202_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_202_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_203_clock; // @[pearray.scala 103:13]
  wire  PE_203_reset; // @[pearray.scala 103:13]
  wire  PE_203_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_203_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_203_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_203_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_203_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_203_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_203_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_203_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_203_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_203_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_203_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_203_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_203_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_204_clock; // @[pearray.scala 103:13]
  wire  PE_204_reset; // @[pearray.scala 103:13]
  wire  PE_204_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_204_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_204_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_204_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_204_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_204_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_204_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_204_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_204_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_204_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_204_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_204_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_204_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_205_clock; // @[pearray.scala 103:13]
  wire  PE_205_reset; // @[pearray.scala 103:13]
  wire  PE_205_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_205_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_205_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_205_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_205_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_205_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_205_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_205_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_205_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_205_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_205_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_205_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_205_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_206_clock; // @[pearray.scala 103:13]
  wire  PE_206_reset; // @[pearray.scala 103:13]
  wire  PE_206_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_206_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_206_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_206_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_206_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_206_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_206_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_206_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_206_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_206_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_206_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_206_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_206_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_207_clock; // @[pearray.scala 103:13]
  wire  PE_207_reset; // @[pearray.scala 103:13]
  wire  PE_207_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_207_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_207_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_207_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_207_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_207_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_207_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_207_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_207_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_207_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_207_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_207_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_207_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_208_clock; // @[pearray.scala 103:13]
  wire  PE_208_reset; // @[pearray.scala 103:13]
  wire  PE_208_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_208_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_208_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_208_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_208_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_208_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_208_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_208_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_208_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_208_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_208_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_208_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_208_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_209_clock; // @[pearray.scala 103:13]
  wire  PE_209_reset; // @[pearray.scala 103:13]
  wire  PE_209_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_209_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_209_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_209_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_209_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_209_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_209_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_209_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_209_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_209_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_209_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_209_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_209_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_210_clock; // @[pearray.scala 103:13]
  wire  PE_210_reset; // @[pearray.scala 103:13]
  wire  PE_210_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_210_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_210_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_210_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_210_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_210_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_210_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_210_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_210_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_210_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_210_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_210_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_210_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_211_clock; // @[pearray.scala 103:13]
  wire  PE_211_reset; // @[pearray.scala 103:13]
  wire  PE_211_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_211_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_211_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_211_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_211_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_211_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_211_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_211_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_211_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_211_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_211_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_211_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_211_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_212_clock; // @[pearray.scala 103:13]
  wire  PE_212_reset; // @[pearray.scala 103:13]
  wire  PE_212_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_212_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_212_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_212_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_212_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_212_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_212_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_212_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_212_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_212_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_212_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_212_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_212_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_213_clock; // @[pearray.scala 103:13]
  wire  PE_213_reset; // @[pearray.scala 103:13]
  wire  PE_213_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_213_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_213_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_213_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_213_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_213_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_213_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_213_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_213_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_213_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_213_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_213_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_213_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_214_clock; // @[pearray.scala 103:13]
  wire  PE_214_reset; // @[pearray.scala 103:13]
  wire  PE_214_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_214_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_214_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_214_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_214_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_214_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_214_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_214_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_214_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_214_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_214_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_214_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_214_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_215_clock; // @[pearray.scala 103:13]
  wire  PE_215_reset; // @[pearray.scala 103:13]
  wire  PE_215_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_215_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_215_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_215_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_215_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_215_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_215_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_215_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_215_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_215_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_215_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_215_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_215_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_216_clock; // @[pearray.scala 103:13]
  wire  PE_216_reset; // @[pearray.scala 103:13]
  wire  PE_216_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_216_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_216_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_216_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_216_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_216_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_216_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_216_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_216_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_216_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_216_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_216_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_216_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_217_clock; // @[pearray.scala 103:13]
  wire  PE_217_reset; // @[pearray.scala 103:13]
  wire  PE_217_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_217_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_217_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_217_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_217_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_217_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_217_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_217_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_217_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_217_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_217_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_217_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_217_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_218_clock; // @[pearray.scala 103:13]
  wire  PE_218_reset; // @[pearray.scala 103:13]
  wire  PE_218_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_218_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_218_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_218_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_218_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_218_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_218_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_218_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_218_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_218_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_218_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_218_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_218_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_219_clock; // @[pearray.scala 103:13]
  wire  PE_219_reset; // @[pearray.scala 103:13]
  wire  PE_219_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_219_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_219_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_219_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_219_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_219_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_219_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_219_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_219_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_219_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_219_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_219_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_219_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_220_clock; // @[pearray.scala 103:13]
  wire  PE_220_reset; // @[pearray.scala 103:13]
  wire  PE_220_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_220_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_220_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_220_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_220_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_220_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_220_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_220_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_220_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_220_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_220_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_220_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_220_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_221_clock; // @[pearray.scala 103:13]
  wire  PE_221_reset; // @[pearray.scala 103:13]
  wire  PE_221_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_221_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_221_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_221_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_221_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_221_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_221_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_221_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_221_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_221_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_221_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_221_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_221_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_222_clock; // @[pearray.scala 103:13]
  wire  PE_222_reset; // @[pearray.scala 103:13]
  wire  PE_222_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_222_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_222_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_222_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_222_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_222_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_222_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_222_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_222_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_222_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_222_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_222_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_222_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_223_clock; // @[pearray.scala 103:13]
  wire  PE_223_reset; // @[pearray.scala 103:13]
  wire  PE_223_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_223_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_223_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_223_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_223_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_223_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_223_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_223_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_223_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_223_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_223_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_223_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_223_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_224_clock; // @[pearray.scala 103:13]
  wire  PE_224_reset; // @[pearray.scala 103:13]
  wire  PE_224_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_224_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_224_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_224_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_224_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_224_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_224_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_224_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_224_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_224_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_224_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_224_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_224_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_225_clock; // @[pearray.scala 103:13]
  wire  PE_225_reset; // @[pearray.scala 103:13]
  wire  PE_225_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_225_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_225_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_225_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_225_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_225_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_225_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_225_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_225_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_225_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_225_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_225_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_225_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_226_clock; // @[pearray.scala 103:13]
  wire  PE_226_reset; // @[pearray.scala 103:13]
  wire  PE_226_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_226_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_226_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_226_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_226_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_226_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_226_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_226_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_226_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_226_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_226_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_226_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_226_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_227_clock; // @[pearray.scala 103:13]
  wire  PE_227_reset; // @[pearray.scala 103:13]
  wire  PE_227_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_227_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_227_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_227_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_227_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_227_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_227_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_227_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_227_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_227_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_227_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_227_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_227_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_228_clock; // @[pearray.scala 103:13]
  wire  PE_228_reset; // @[pearray.scala 103:13]
  wire  PE_228_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_228_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_228_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_228_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_228_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_228_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_228_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_228_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_228_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_228_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_228_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_228_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_228_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_229_clock; // @[pearray.scala 103:13]
  wire  PE_229_reset; // @[pearray.scala 103:13]
  wire  PE_229_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_229_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_229_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_229_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_229_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_229_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_229_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_229_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_229_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_229_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_229_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_229_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_229_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_230_clock; // @[pearray.scala 103:13]
  wire  PE_230_reset; // @[pearray.scala 103:13]
  wire  PE_230_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_230_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_230_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_230_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_230_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_230_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_230_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_230_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_230_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_230_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_230_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_230_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_230_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_231_clock; // @[pearray.scala 103:13]
  wire  PE_231_reset; // @[pearray.scala 103:13]
  wire  PE_231_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_231_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_231_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_231_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_231_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_231_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_231_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_231_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_231_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_231_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_231_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_231_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_231_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_232_clock; // @[pearray.scala 103:13]
  wire  PE_232_reset; // @[pearray.scala 103:13]
  wire  PE_232_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_232_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_232_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_232_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_232_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_232_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_232_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_232_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_232_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_232_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_232_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_232_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_232_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_233_clock; // @[pearray.scala 103:13]
  wire  PE_233_reset; // @[pearray.scala 103:13]
  wire  PE_233_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_233_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_233_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_233_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_233_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_233_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_233_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_233_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_233_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_233_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_233_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_233_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_233_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_234_clock; // @[pearray.scala 103:13]
  wire  PE_234_reset; // @[pearray.scala 103:13]
  wire  PE_234_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_234_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_234_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_234_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_234_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_234_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_234_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_234_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_234_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_234_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_234_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_234_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_234_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_235_clock; // @[pearray.scala 103:13]
  wire  PE_235_reset; // @[pearray.scala 103:13]
  wire  PE_235_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_235_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_235_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_235_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_235_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_235_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_235_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_235_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_235_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_235_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_235_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_235_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_235_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_236_clock; // @[pearray.scala 103:13]
  wire  PE_236_reset; // @[pearray.scala 103:13]
  wire  PE_236_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_236_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_236_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_236_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_236_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_236_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_236_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_236_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_236_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_236_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_236_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_236_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_236_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_237_clock; // @[pearray.scala 103:13]
  wire  PE_237_reset; // @[pearray.scala 103:13]
  wire  PE_237_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_237_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_237_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_237_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_237_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_237_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_237_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_237_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_237_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_237_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_237_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_237_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_237_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_238_clock; // @[pearray.scala 103:13]
  wire  PE_238_reset; // @[pearray.scala 103:13]
  wire  PE_238_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_238_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_238_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_238_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_238_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_238_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_238_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_238_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_238_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_238_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_238_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_238_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_238_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_239_clock; // @[pearray.scala 103:13]
  wire  PE_239_reset; // @[pearray.scala 103:13]
  wire  PE_239_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_239_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_239_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_239_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_239_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_239_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_239_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_239_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_239_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_239_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_239_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_239_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_239_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_240_clock; // @[pearray.scala 103:13]
  wire  PE_240_reset; // @[pearray.scala 103:13]
  wire  PE_240_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_240_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_240_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_240_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_240_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_240_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_240_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_240_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_240_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_240_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_240_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_240_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_240_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_241_clock; // @[pearray.scala 103:13]
  wire  PE_241_reset; // @[pearray.scala 103:13]
  wire  PE_241_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_241_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_241_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_241_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_241_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_241_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_241_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_241_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_241_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_241_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_241_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_241_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_241_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_242_clock; // @[pearray.scala 103:13]
  wire  PE_242_reset; // @[pearray.scala 103:13]
  wire  PE_242_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_242_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_242_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_242_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_242_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_242_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_242_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_242_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_242_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_242_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_242_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_242_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_242_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_243_clock; // @[pearray.scala 103:13]
  wire  PE_243_reset; // @[pearray.scala 103:13]
  wire  PE_243_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_243_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_243_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_243_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_243_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_243_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_243_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_243_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_243_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_243_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_243_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_243_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_243_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_244_clock; // @[pearray.scala 103:13]
  wire  PE_244_reset; // @[pearray.scala 103:13]
  wire  PE_244_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_244_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_244_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_244_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_244_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_244_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_244_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_244_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_244_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_244_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_244_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_244_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_244_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_245_clock; // @[pearray.scala 103:13]
  wire  PE_245_reset; // @[pearray.scala 103:13]
  wire  PE_245_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_245_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_245_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_245_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_245_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_245_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_245_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_245_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_245_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_245_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_245_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_245_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_245_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_246_clock; // @[pearray.scala 103:13]
  wire  PE_246_reset; // @[pearray.scala 103:13]
  wire  PE_246_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_246_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_246_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_246_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_246_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_246_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_246_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_246_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_246_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_246_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_246_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_246_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_246_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_247_clock; // @[pearray.scala 103:13]
  wire  PE_247_reset; // @[pearray.scala 103:13]
  wire  PE_247_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_247_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_247_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_247_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_247_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_247_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_247_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_247_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_247_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_247_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_247_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_247_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_247_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_248_clock; // @[pearray.scala 103:13]
  wire  PE_248_reset; // @[pearray.scala 103:13]
  wire  PE_248_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_248_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_248_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_248_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_248_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_248_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_248_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_248_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_248_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_248_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_248_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_248_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_248_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_249_clock; // @[pearray.scala 103:13]
  wire  PE_249_reset; // @[pearray.scala 103:13]
  wire  PE_249_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_249_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_249_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_249_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_249_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_249_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_249_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_249_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_249_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_249_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_249_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_249_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_249_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_250_clock; // @[pearray.scala 103:13]
  wire  PE_250_reset; // @[pearray.scala 103:13]
  wire  PE_250_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_250_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_250_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_250_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_250_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_250_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_250_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_250_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_250_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_250_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_250_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_250_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_250_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_251_clock; // @[pearray.scala 103:13]
  wire  PE_251_reset; // @[pearray.scala 103:13]
  wire  PE_251_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_251_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_251_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_251_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_251_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_251_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_251_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_251_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_251_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_251_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_251_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_251_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_251_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_252_clock; // @[pearray.scala 103:13]
  wire  PE_252_reset; // @[pearray.scala 103:13]
  wire  PE_252_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_252_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_252_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_252_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_252_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_252_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_252_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_252_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_252_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_252_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_252_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_252_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_252_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_253_clock; // @[pearray.scala 103:13]
  wire  PE_253_reset; // @[pearray.scala 103:13]
  wire  PE_253_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_253_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_253_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_253_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_253_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_253_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_253_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_253_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_253_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_253_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_253_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_253_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_253_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_254_clock; // @[pearray.scala 103:13]
  wire  PE_254_reset; // @[pearray.scala 103:13]
  wire  PE_254_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_254_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_254_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_254_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_254_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_254_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_254_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_254_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_254_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_254_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_254_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_254_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_254_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_255_clock; // @[pearray.scala 103:13]
  wire  PE_255_reset; // @[pearray.scala 103:13]
  wire  PE_255_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_255_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_255_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_255_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_255_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_255_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_255_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_255_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_255_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_255_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_255_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_255_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_255_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PENetwork_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_15_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_15_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_24_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_24_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_25_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_25_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_26_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_26_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_27_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_27_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_28_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_28_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_29_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_29_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_30_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_30_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_31_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_31_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_32_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_32_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_33_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_33_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_34_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_34_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_35_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_35_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_36_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_36_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_37_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_37_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_38_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_38_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_39_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_39_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_40_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_40_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_41_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_41_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_42_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_42_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_43_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_43_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_44_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_44_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_45_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_45_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_46_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_46_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_8_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_8_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_8_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_8_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_9_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_9_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_9_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_9_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_10_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_10_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_10_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_10_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_11_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_11_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_11_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_11_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_12_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_12_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_12_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_12_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_13_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_13_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_13_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_13_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_14_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_14_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_14_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_14_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_pes_15_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_pes_15_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_47_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_47_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  MemController_clock; // @[pearray.scala 212:15]
  wire  MemController_reset; // @[pearray.scala 212:15]
  wire  MemController_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_1_clock; // @[pearray.scala 212:15]
  wire  MemController_1_reset; // @[pearray.scala 212:15]
  wire  MemController_1_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_1_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_1_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_1_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_1_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_1_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_2_clock; // @[pearray.scala 212:15]
  wire  MemController_2_reset; // @[pearray.scala 212:15]
  wire  MemController_2_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_2_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_2_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_2_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_2_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_2_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_3_clock; // @[pearray.scala 212:15]
  wire  MemController_3_reset; // @[pearray.scala 212:15]
  wire  MemController_3_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_3_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_3_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_3_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_3_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_3_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_4_clock; // @[pearray.scala 212:15]
  wire  MemController_4_reset; // @[pearray.scala 212:15]
  wire  MemController_4_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_4_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_4_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_4_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_4_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_4_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_5_clock; // @[pearray.scala 212:15]
  wire  MemController_5_reset; // @[pearray.scala 212:15]
  wire  MemController_5_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_5_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_5_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_5_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_5_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_5_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_6_clock; // @[pearray.scala 212:15]
  wire  MemController_6_reset; // @[pearray.scala 212:15]
  wire  MemController_6_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_6_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_6_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_6_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_6_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_6_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_7_clock; // @[pearray.scala 212:15]
  wire  MemController_7_reset; // @[pearray.scala 212:15]
  wire  MemController_7_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_7_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_7_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_7_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_7_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_7_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_8_clock; // @[pearray.scala 212:15]
  wire  MemController_8_reset; // @[pearray.scala 212:15]
  wire  MemController_8_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_8_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_8_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_8_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_8_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_8_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_9_clock; // @[pearray.scala 212:15]
  wire  MemController_9_reset; // @[pearray.scala 212:15]
  wire  MemController_9_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_9_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_9_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_9_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_9_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_9_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_10_clock; // @[pearray.scala 212:15]
  wire  MemController_10_reset; // @[pearray.scala 212:15]
  wire  MemController_10_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_10_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_10_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_10_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_10_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_10_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_11_clock; // @[pearray.scala 212:15]
  wire  MemController_11_reset; // @[pearray.scala 212:15]
  wire  MemController_11_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_11_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_11_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_11_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_11_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_11_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_12_clock; // @[pearray.scala 212:15]
  wire  MemController_12_reset; // @[pearray.scala 212:15]
  wire  MemController_12_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_12_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_12_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_12_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_12_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_12_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_13_clock; // @[pearray.scala 212:15]
  wire  MemController_13_reset; // @[pearray.scala 212:15]
  wire  MemController_13_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_13_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_13_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_13_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_13_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_13_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_14_clock; // @[pearray.scala 212:15]
  wire  MemController_14_reset; // @[pearray.scala 212:15]
  wire  MemController_14_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_14_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_14_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_14_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_14_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_14_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_15_clock; // @[pearray.scala 212:15]
  wire  MemController_15_reset; // @[pearray.scala 212:15]
  wire  MemController_15_io_rd_valid; // @[pearray.scala 212:15]
  wire  MemController_15_io_wr_valid; // @[pearray.scala 212:15]
  wire  MemController_15_io_rd_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_15_io_rd_data_bits; // @[pearray.scala 212:15]
  wire  MemController_15_io_wr_data_valid; // @[pearray.scala 212:15]
  wire [15:0] MemController_15_io_wr_data_bits; // @[pearray.scala 212:15]
  wire  MemController_16_clock; // @[pearray.scala 210:15]
  wire  MemController_16_reset; // @[pearray.scala 210:15]
  wire  MemController_16_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_16_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_16_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_16_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_16_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_16_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_17_clock; // @[pearray.scala 210:15]
  wire  MemController_17_reset; // @[pearray.scala 210:15]
  wire  MemController_17_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_17_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_17_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_17_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_17_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_17_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_18_clock; // @[pearray.scala 210:15]
  wire  MemController_18_reset; // @[pearray.scala 210:15]
  wire  MemController_18_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_18_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_18_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_18_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_18_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_18_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_19_clock; // @[pearray.scala 210:15]
  wire  MemController_19_reset; // @[pearray.scala 210:15]
  wire  MemController_19_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_19_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_19_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_19_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_19_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_19_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_20_clock; // @[pearray.scala 210:15]
  wire  MemController_20_reset; // @[pearray.scala 210:15]
  wire  MemController_20_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_20_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_20_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_20_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_20_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_20_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_21_clock; // @[pearray.scala 210:15]
  wire  MemController_21_reset; // @[pearray.scala 210:15]
  wire  MemController_21_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_21_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_21_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_21_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_21_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_21_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_22_clock; // @[pearray.scala 210:15]
  wire  MemController_22_reset; // @[pearray.scala 210:15]
  wire  MemController_22_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_22_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_22_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_22_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_22_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_22_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_23_clock; // @[pearray.scala 210:15]
  wire  MemController_23_reset; // @[pearray.scala 210:15]
  wire  MemController_23_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_23_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_23_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_23_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_23_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_23_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_24_clock; // @[pearray.scala 210:15]
  wire  MemController_24_reset; // @[pearray.scala 210:15]
  wire  MemController_24_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_24_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_24_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_24_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_24_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_24_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_25_clock; // @[pearray.scala 210:15]
  wire  MemController_25_reset; // @[pearray.scala 210:15]
  wire  MemController_25_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_25_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_25_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_25_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_25_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_25_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_26_clock; // @[pearray.scala 210:15]
  wire  MemController_26_reset; // @[pearray.scala 210:15]
  wire  MemController_26_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_26_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_26_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_26_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_26_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_26_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_27_clock; // @[pearray.scala 210:15]
  wire  MemController_27_reset; // @[pearray.scala 210:15]
  wire  MemController_27_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_27_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_27_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_27_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_27_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_27_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_28_clock; // @[pearray.scala 210:15]
  wire  MemController_28_reset; // @[pearray.scala 210:15]
  wire  MemController_28_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_28_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_28_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_28_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_28_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_28_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_29_clock; // @[pearray.scala 210:15]
  wire  MemController_29_reset; // @[pearray.scala 210:15]
  wire  MemController_29_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_29_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_29_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_29_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_29_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_29_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_30_clock; // @[pearray.scala 210:15]
  wire  MemController_30_reset; // @[pearray.scala 210:15]
  wire  MemController_30_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_30_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_30_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_30_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_30_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_30_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_31_clock; // @[pearray.scala 210:15]
  wire  MemController_31_reset; // @[pearray.scala 210:15]
  wire  MemController_31_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_31_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_31_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_31_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_31_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_31_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_32_clock; // @[pearray.scala 210:15]
  wire  MemController_32_reset; // @[pearray.scala 210:15]
  wire  MemController_32_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_32_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_32_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_32_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_32_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_32_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_33_clock; // @[pearray.scala 210:15]
  wire  MemController_33_reset; // @[pearray.scala 210:15]
  wire  MemController_33_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_33_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_33_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_33_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_33_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_33_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_34_clock; // @[pearray.scala 210:15]
  wire  MemController_34_reset; // @[pearray.scala 210:15]
  wire  MemController_34_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_34_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_34_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_34_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_34_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_34_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_35_clock; // @[pearray.scala 210:15]
  wire  MemController_35_reset; // @[pearray.scala 210:15]
  wire  MemController_35_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_35_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_35_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_35_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_35_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_35_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_36_clock; // @[pearray.scala 210:15]
  wire  MemController_36_reset; // @[pearray.scala 210:15]
  wire  MemController_36_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_36_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_36_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_36_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_36_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_36_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_37_clock; // @[pearray.scala 210:15]
  wire  MemController_37_reset; // @[pearray.scala 210:15]
  wire  MemController_37_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_37_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_37_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_37_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_37_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_37_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_38_clock; // @[pearray.scala 210:15]
  wire  MemController_38_reset; // @[pearray.scala 210:15]
  wire  MemController_38_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_38_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_38_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_38_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_38_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_38_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_39_clock; // @[pearray.scala 210:15]
  wire  MemController_39_reset; // @[pearray.scala 210:15]
  wire  MemController_39_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_39_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_39_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_39_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_39_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_39_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_40_clock; // @[pearray.scala 210:15]
  wire  MemController_40_reset; // @[pearray.scala 210:15]
  wire  MemController_40_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_40_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_40_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_40_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_40_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_40_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_41_clock; // @[pearray.scala 210:15]
  wire  MemController_41_reset; // @[pearray.scala 210:15]
  wire  MemController_41_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_41_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_41_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_41_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_41_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_41_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_42_clock; // @[pearray.scala 210:15]
  wire  MemController_42_reset; // @[pearray.scala 210:15]
  wire  MemController_42_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_42_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_42_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_42_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_42_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_42_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_43_clock; // @[pearray.scala 210:15]
  wire  MemController_43_reset; // @[pearray.scala 210:15]
  wire  MemController_43_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_43_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_43_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_43_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_43_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_43_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_44_clock; // @[pearray.scala 210:15]
  wire  MemController_44_reset; // @[pearray.scala 210:15]
  wire  MemController_44_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_44_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_44_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_44_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_44_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_44_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_45_clock; // @[pearray.scala 210:15]
  wire  MemController_45_reset; // @[pearray.scala 210:15]
  wire  MemController_45_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_45_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_45_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_45_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_45_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_45_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_46_clock; // @[pearray.scala 210:15]
  wire  MemController_46_reset; // @[pearray.scala 210:15]
  wire  MemController_46_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_46_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_46_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_46_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_46_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_46_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  MemController_47_clock; // @[pearray.scala 210:15]
  wire  MemController_47_reset; // @[pearray.scala 210:15]
  wire  MemController_47_io_rd_valid; // @[pearray.scala 210:15]
  wire  MemController_47_io_wr_valid; // @[pearray.scala 210:15]
  wire  MemController_47_io_rd_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_47_io_rd_data_bits; // @[pearray.scala 210:15]
  wire  MemController_47_io_wr_data_valid; // @[pearray.scala 210:15]
  wire [15:0] MemController_47_io_wr_data_bits; // @[pearray.scala 210:15]
  wire  _T_3 = MultiDimTime_io_index_1 == 18'h0; // @[pearray.scala 182:41]
  wire  _T_4 = MultiDimTime_io_index_0 == 18'h0; // @[pearray.scala 182:89]
  wire  _T_5 = _T_3 & _T_4; // @[pearray.scala 182:67]
  reg  _T_12_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_0;
  reg  _T_12_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1;
  reg  _T_12_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_2;
  reg  _T_12_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_3;
  wire  _T_13 = MultiDimTime_io_index_1 == 18'h1; // @[pearray.scala 182:41]
  wire  _T_15 = _T_13 & _T_4; // @[pearray.scala 182:67]
  reg  _T_22_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_4;
  reg  _T_22_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_5;
  reg  _T_22_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_6;
  reg  _T_22_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_7;
  wire  _T_23 = MultiDimTime_io_index_1 == 18'h2; // @[pearray.scala 182:41]
  wire  _T_25 = _T_23 & _T_4; // @[pearray.scala 182:67]
  reg  _T_32_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_8;
  reg  _T_32_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_9;
  reg  _T_32_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_10;
  reg  _T_32_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_11;
  wire  _T_33 = MultiDimTime_io_index_1 == 18'h3; // @[pearray.scala 182:41]
  wire  _T_35 = _T_33 & _T_4; // @[pearray.scala 182:67]
  reg  _T_42_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_12;
  reg  _T_42_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_13;
  reg  _T_42_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_14;
  reg  _T_42_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_15;
  wire  _T_43 = MultiDimTime_io_index_1 == 18'h4; // @[pearray.scala 182:41]
  wire  _T_45 = _T_43 & _T_4; // @[pearray.scala 182:67]
  reg  _T_52_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_16;
  reg  _T_52_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_17;
  reg  _T_52_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_18;
  reg  _T_52_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_19;
  wire  _T_53 = MultiDimTime_io_index_1 == 18'h5; // @[pearray.scala 182:41]
  wire  _T_55 = _T_53 & _T_4; // @[pearray.scala 182:67]
  reg  _T_62_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_20;
  reg  _T_62_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_21;
  reg  _T_62_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_22;
  reg  _T_62_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_23;
  wire  _T_63 = MultiDimTime_io_index_1 == 18'h6; // @[pearray.scala 182:41]
  wire  _T_65 = _T_63 & _T_4; // @[pearray.scala 182:67]
  reg  _T_72_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_24;
  reg  _T_72_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_25;
  reg  _T_72_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_26;
  reg  _T_72_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_27;
  wire  _T_73 = MultiDimTime_io_index_1 == 18'h7; // @[pearray.scala 182:41]
  wire  _T_75 = _T_73 & _T_4; // @[pearray.scala 182:67]
  reg  _T_82_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_28;
  reg  _T_82_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_29;
  reg  _T_82_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_30;
  reg  _T_82_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_31;
  wire  _T_83 = MultiDimTime_io_index_1 == 18'h8; // @[pearray.scala 182:41]
  wire  _T_85 = _T_83 & _T_4; // @[pearray.scala 182:67]
  reg  _T_92_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_32;
  reg  _T_92_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_33;
  reg  _T_92_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_34;
  reg  _T_92_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_35;
  wire  _T_93 = MultiDimTime_io_index_1 == 18'h9; // @[pearray.scala 182:41]
  wire  _T_95 = _T_93 & _T_4; // @[pearray.scala 182:67]
  reg  _T_102_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_36;
  reg  _T_102_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_37;
  reg  _T_102_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_38;
  reg  _T_102_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_39;
  wire  _T_103 = MultiDimTime_io_index_1 == 18'ha; // @[pearray.scala 182:41]
  wire  _T_105 = _T_103 & _T_4; // @[pearray.scala 182:67]
  reg  _T_112_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_40;
  reg  _T_112_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_41;
  reg  _T_112_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_42;
  reg  _T_112_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_43;
  wire  _T_113 = MultiDimTime_io_index_1 == 18'hb; // @[pearray.scala 182:41]
  wire  _T_115 = _T_113 & _T_4; // @[pearray.scala 182:67]
  reg  _T_122_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_44;
  reg  _T_122_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_45;
  reg  _T_122_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_46;
  reg  _T_122_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_47;
  wire  _T_123 = MultiDimTime_io_index_1 == 18'hc; // @[pearray.scala 182:41]
  wire  _T_125 = _T_123 & _T_4; // @[pearray.scala 182:67]
  reg  _T_132_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_48;
  reg  _T_132_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_49;
  reg  _T_132_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_50;
  reg  _T_132_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_51;
  wire  _T_133 = MultiDimTime_io_index_1 == 18'hd; // @[pearray.scala 182:41]
  wire  _T_135 = _T_133 & _T_4; // @[pearray.scala 182:67]
  reg  _T_142_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_52;
  reg  _T_142_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_53;
  reg  _T_142_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_54;
  reg  _T_142_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_55;
  wire  _T_143 = MultiDimTime_io_index_1 == 18'he; // @[pearray.scala 182:41]
  wire  _T_145 = _T_143 & _T_4; // @[pearray.scala 182:67]
  reg  _T_152_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_56;
  reg  _T_152_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_57;
  reg  _T_152_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_58;
  reg  _T_152_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_59;
  wire  _T_153 = MultiDimTime_io_index_1 == 18'hf; // @[pearray.scala 182:41]
  wire  _T_155 = _T_153 & _T_4; // @[pearray.scala 182:67]
  reg  _T_162_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_60;
  reg  _T_162_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_61;
  reg  _T_162_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_62;
  reg  _T_162_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_63;
  reg  _T_172_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_64;
  reg  _T_172_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_65;
  reg  _T_172_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_66;
  reg  _T_172_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_67;
  reg  _T_182_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_68;
  reg  _T_182_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_69;
  reg  _T_182_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_70;
  reg  _T_182_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_71;
  reg  _T_192_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_72;
  reg  _T_192_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_73;
  reg  _T_192_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_74;
  reg  _T_192_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_75;
  reg  _T_202_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_76;
  reg  _T_202_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_77;
  reg  _T_202_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_78;
  reg  _T_202_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_79;
  reg  _T_212_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_80;
  reg  _T_212_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_81;
  reg  _T_212_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_82;
  reg  _T_212_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_83;
  reg  _T_222_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_84;
  reg  _T_222_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_85;
  reg  _T_222_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_86;
  reg  _T_222_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_87;
  reg  _T_232_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_88;
  reg  _T_232_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_89;
  reg  _T_232_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_90;
  reg  _T_232_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_91;
  reg  _T_242_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_92;
  reg  _T_242_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_93;
  reg  _T_242_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_94;
  reg  _T_242_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_95;
  reg  _T_252_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_96;
  reg  _T_252_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_97;
  reg  _T_252_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_98;
  reg  _T_252_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_99;
  reg  _T_262_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_100;
  reg  _T_262_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_101;
  reg  _T_262_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_102;
  reg  _T_262_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_103;
  reg  _T_272_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_104;
  reg  _T_272_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_105;
  reg  _T_272_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_106;
  reg  _T_272_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_107;
  reg  _T_282_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_108;
  reg  _T_282_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_109;
  reg  _T_282_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_110;
  reg  _T_282_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_111;
  reg  _T_292_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_112;
  reg  _T_292_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_113;
  reg  _T_292_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_114;
  reg  _T_292_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_115;
  reg  _T_302_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_116;
  reg  _T_302_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_117;
  reg  _T_302_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_118;
  reg  _T_302_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_119;
  reg  _T_312_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_120;
  reg  _T_312_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_121;
  reg  _T_312_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_122;
  reg  _T_312_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_123;
  wire  _T_313 = MultiDimTime_io_index_1 == 18'h10; // @[pearray.scala 182:41]
  wire  _T_315 = _T_313 & _T_4; // @[pearray.scala 182:67]
  reg  _T_322_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_124;
  reg  _T_322_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_125;
  reg  _T_322_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_126;
  reg  _T_322_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_127;
  reg  _T_332_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_128;
  reg  _T_332_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_129;
  reg  _T_332_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_130;
  reg  _T_332_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_131;
  reg  _T_342_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_132;
  reg  _T_342_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_133;
  reg  _T_342_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_134;
  reg  _T_342_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_135;
  reg  _T_352_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_136;
  reg  _T_352_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_137;
  reg  _T_352_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_138;
  reg  _T_352_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_139;
  reg  _T_362_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_140;
  reg  _T_362_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_141;
  reg  _T_362_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_142;
  reg  _T_362_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_143;
  reg  _T_372_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_144;
  reg  _T_372_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_145;
  reg  _T_372_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_146;
  reg  _T_372_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_147;
  reg  _T_382_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_148;
  reg  _T_382_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_149;
  reg  _T_382_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_150;
  reg  _T_382_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_151;
  reg  _T_392_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_152;
  reg  _T_392_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_153;
  reg  _T_392_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_154;
  reg  _T_392_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_155;
  reg  _T_402_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_156;
  reg  _T_402_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_157;
  reg  _T_402_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_158;
  reg  _T_402_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_159;
  reg  _T_412_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_160;
  reg  _T_412_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_161;
  reg  _T_412_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_162;
  reg  _T_412_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_163;
  reg  _T_422_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_164;
  reg  _T_422_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_165;
  reg  _T_422_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_166;
  reg  _T_422_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_167;
  reg  _T_432_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_168;
  reg  _T_432_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_169;
  reg  _T_432_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_170;
  reg  _T_432_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_171;
  reg  _T_442_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_172;
  reg  _T_442_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_173;
  reg  _T_442_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_174;
  reg  _T_442_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_175;
  reg  _T_452_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_176;
  reg  _T_452_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_177;
  reg  _T_452_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_178;
  reg  _T_452_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_179;
  reg  _T_462_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_180;
  reg  _T_462_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_181;
  reg  _T_462_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_182;
  reg  _T_462_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_183;
  reg  _T_472_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_184;
  reg  _T_472_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_185;
  reg  _T_472_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_186;
  reg  _T_472_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_187;
  wire  _T_473 = MultiDimTime_io_index_1 == 18'h11; // @[pearray.scala 182:41]
  wire  _T_475 = _T_473 & _T_4; // @[pearray.scala 182:67]
  reg  _T_482_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_188;
  reg  _T_482_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_189;
  reg  _T_482_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_190;
  reg  _T_482_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_191;
  reg  _T_492_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_192;
  reg  _T_492_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_193;
  reg  _T_492_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_194;
  reg  _T_492_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_195;
  reg  _T_502_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_196;
  reg  _T_502_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_197;
  reg  _T_502_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_198;
  reg  _T_502_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_199;
  reg  _T_512_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_200;
  reg  _T_512_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_201;
  reg  _T_512_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_202;
  reg  _T_512_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_203;
  reg  _T_522_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_204;
  reg  _T_522_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_205;
  reg  _T_522_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_206;
  reg  _T_522_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_207;
  reg  _T_532_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_208;
  reg  _T_532_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_209;
  reg  _T_532_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_210;
  reg  _T_532_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_211;
  reg  _T_542_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_212;
  reg  _T_542_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_213;
  reg  _T_542_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_214;
  reg  _T_542_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_215;
  reg  _T_552_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_216;
  reg  _T_552_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_217;
  reg  _T_552_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_218;
  reg  _T_552_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_219;
  reg  _T_562_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_220;
  reg  _T_562_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_221;
  reg  _T_562_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_222;
  reg  _T_562_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_223;
  reg  _T_572_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_224;
  reg  _T_572_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_225;
  reg  _T_572_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_226;
  reg  _T_572_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_227;
  reg  _T_582_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_228;
  reg  _T_582_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_229;
  reg  _T_582_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_230;
  reg  _T_582_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_231;
  reg  _T_592_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_232;
  reg  _T_592_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_233;
  reg  _T_592_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_234;
  reg  _T_592_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_235;
  reg  _T_602_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_236;
  reg  _T_602_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_237;
  reg  _T_602_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_238;
  reg  _T_602_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_239;
  reg  _T_612_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_240;
  reg  _T_612_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_241;
  reg  _T_612_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_242;
  reg  _T_612_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_243;
  reg  _T_622_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_244;
  reg  _T_622_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_245;
  reg  _T_622_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_246;
  reg  _T_622_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_247;
  reg  _T_632_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_248;
  reg  _T_632_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_249;
  reg  _T_632_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_250;
  reg  _T_632_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_251;
  wire  _T_633 = MultiDimTime_io_index_1 == 18'h12; // @[pearray.scala 182:41]
  wire  _T_635 = _T_633 & _T_4; // @[pearray.scala 182:67]
  reg  _T_642_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_252;
  reg  _T_642_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_253;
  reg  _T_642_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_254;
  reg  _T_642_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_255;
  reg  _T_652_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_256;
  reg  _T_652_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_257;
  reg  _T_652_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_258;
  reg  _T_652_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_259;
  reg  _T_662_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_260;
  reg  _T_662_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_261;
  reg  _T_662_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_262;
  reg  _T_662_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_263;
  reg  _T_672_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_264;
  reg  _T_672_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_265;
  reg  _T_672_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_266;
  reg  _T_672_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_267;
  reg  _T_682_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_268;
  reg  _T_682_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_269;
  reg  _T_682_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_270;
  reg  _T_682_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_271;
  reg  _T_692_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_272;
  reg  _T_692_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_273;
  reg  _T_692_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_274;
  reg  _T_692_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_275;
  reg  _T_702_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_276;
  reg  _T_702_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_277;
  reg  _T_702_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_278;
  reg  _T_702_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_279;
  reg  _T_712_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_280;
  reg  _T_712_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_281;
  reg  _T_712_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_282;
  reg  _T_712_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_283;
  reg  _T_722_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_284;
  reg  _T_722_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_285;
  reg  _T_722_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_286;
  reg  _T_722_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_287;
  reg  _T_732_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_288;
  reg  _T_732_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_289;
  reg  _T_732_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_290;
  reg  _T_732_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_291;
  reg  _T_742_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_292;
  reg  _T_742_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_293;
  reg  _T_742_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_294;
  reg  _T_742_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_295;
  reg  _T_752_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_296;
  reg  _T_752_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_297;
  reg  _T_752_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_298;
  reg  _T_752_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_299;
  reg  _T_762_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_300;
  reg  _T_762_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_301;
  reg  _T_762_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_302;
  reg  _T_762_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_303;
  reg  _T_772_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_304;
  reg  _T_772_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_305;
  reg  _T_772_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_306;
  reg  _T_772_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_307;
  reg  _T_782_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_308;
  reg  _T_782_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_309;
  reg  _T_782_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_310;
  reg  _T_782_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_311;
  reg  _T_792_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_312;
  reg  _T_792_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_313;
  reg  _T_792_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_314;
  reg  _T_792_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_315;
  wire  _T_793 = MultiDimTime_io_index_1 == 18'h13; // @[pearray.scala 182:41]
  wire  _T_795 = _T_793 & _T_4; // @[pearray.scala 182:67]
  reg  _T_802_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_316;
  reg  _T_802_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_317;
  reg  _T_802_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_318;
  reg  _T_802_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_319;
  reg  _T_812_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_320;
  reg  _T_812_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_321;
  reg  _T_812_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_322;
  reg  _T_812_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_323;
  reg  _T_822_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_324;
  reg  _T_822_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_325;
  reg  _T_822_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_326;
  reg  _T_822_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_327;
  reg  _T_832_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_328;
  reg  _T_832_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_329;
  reg  _T_832_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_330;
  reg  _T_832_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_331;
  reg  _T_842_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_332;
  reg  _T_842_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_333;
  reg  _T_842_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_334;
  reg  _T_842_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_335;
  reg  _T_852_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_336;
  reg  _T_852_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_337;
  reg  _T_852_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_338;
  reg  _T_852_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_339;
  reg  _T_862_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_340;
  reg  _T_862_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_341;
  reg  _T_862_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_342;
  reg  _T_862_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_343;
  reg  _T_872_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_344;
  reg  _T_872_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_345;
  reg  _T_872_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_346;
  reg  _T_872_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_347;
  reg  _T_882_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_348;
  reg  _T_882_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_349;
  reg  _T_882_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_350;
  reg  _T_882_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_351;
  reg  _T_892_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_352;
  reg  _T_892_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_353;
  reg  _T_892_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_354;
  reg  _T_892_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_355;
  reg  _T_902_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_356;
  reg  _T_902_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_357;
  reg  _T_902_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_358;
  reg  _T_902_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_359;
  reg  _T_912_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_360;
  reg  _T_912_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_361;
  reg  _T_912_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_362;
  reg  _T_912_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_363;
  reg  _T_922_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_364;
  reg  _T_922_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_365;
  reg  _T_922_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_366;
  reg  _T_922_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_367;
  reg  _T_932_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_368;
  reg  _T_932_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_369;
  reg  _T_932_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_370;
  reg  _T_932_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_371;
  reg  _T_942_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_372;
  reg  _T_942_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_373;
  reg  _T_942_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_374;
  reg  _T_942_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_375;
  reg  _T_952_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_376;
  reg  _T_952_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_377;
  reg  _T_952_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_378;
  reg  _T_952_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_379;
  wire  _T_953 = MultiDimTime_io_index_1 == 18'h14; // @[pearray.scala 182:41]
  wire  _T_955 = _T_953 & _T_4; // @[pearray.scala 182:67]
  reg  _T_962_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_380;
  reg  _T_962_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_381;
  reg  _T_962_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_382;
  reg  _T_962_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_383;
  reg  _T_972_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_384;
  reg  _T_972_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_385;
  reg  _T_972_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_386;
  reg  _T_972_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_387;
  reg  _T_982_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_388;
  reg  _T_982_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_389;
  reg  _T_982_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_390;
  reg  _T_982_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_391;
  reg  _T_992_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_392;
  reg  _T_992_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_393;
  reg  _T_992_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_394;
  reg  _T_992_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_395;
  reg  _T_1002_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_396;
  reg  _T_1002_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_397;
  reg  _T_1002_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_398;
  reg  _T_1002_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_399;
  reg  _T_1012_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_400;
  reg  _T_1012_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_401;
  reg  _T_1012_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_402;
  reg  _T_1012_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_403;
  reg  _T_1022_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_404;
  reg  _T_1022_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_405;
  reg  _T_1022_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_406;
  reg  _T_1022_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_407;
  reg  _T_1032_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_408;
  reg  _T_1032_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_409;
  reg  _T_1032_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_410;
  reg  _T_1032_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_411;
  reg  _T_1042_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_412;
  reg  _T_1042_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_413;
  reg  _T_1042_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_414;
  reg  _T_1042_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_415;
  reg  _T_1052_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_416;
  reg  _T_1052_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_417;
  reg  _T_1052_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_418;
  reg  _T_1052_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_419;
  reg  _T_1062_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_420;
  reg  _T_1062_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_421;
  reg  _T_1062_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_422;
  reg  _T_1062_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_423;
  reg  _T_1072_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_424;
  reg  _T_1072_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_425;
  reg  _T_1072_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_426;
  reg  _T_1072_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_427;
  reg  _T_1082_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_428;
  reg  _T_1082_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_429;
  reg  _T_1082_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_430;
  reg  _T_1082_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_431;
  reg  _T_1092_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_432;
  reg  _T_1092_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_433;
  reg  _T_1092_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_434;
  reg  _T_1092_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_435;
  reg  _T_1102_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_436;
  reg  _T_1102_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_437;
  reg  _T_1102_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_438;
  reg  _T_1102_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_439;
  reg  _T_1112_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_440;
  reg  _T_1112_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_441;
  reg  _T_1112_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_442;
  reg  _T_1112_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_443;
  wire  _T_1113 = MultiDimTime_io_index_1 == 18'h15; // @[pearray.scala 182:41]
  wire  _T_1115 = _T_1113 & _T_4; // @[pearray.scala 182:67]
  reg  _T_1122_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_444;
  reg  _T_1122_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_445;
  reg  _T_1122_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_446;
  reg  _T_1122_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_447;
  reg  _T_1132_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_448;
  reg  _T_1132_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_449;
  reg  _T_1132_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_450;
  reg  _T_1132_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_451;
  reg  _T_1142_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_452;
  reg  _T_1142_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_453;
  reg  _T_1142_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_454;
  reg  _T_1142_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_455;
  reg  _T_1152_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_456;
  reg  _T_1152_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_457;
  reg  _T_1152_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_458;
  reg  _T_1152_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_459;
  reg  _T_1162_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_460;
  reg  _T_1162_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_461;
  reg  _T_1162_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_462;
  reg  _T_1162_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_463;
  reg  _T_1172_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_464;
  reg  _T_1172_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_465;
  reg  _T_1172_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_466;
  reg  _T_1172_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_467;
  reg  _T_1182_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_468;
  reg  _T_1182_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_469;
  reg  _T_1182_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_470;
  reg  _T_1182_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_471;
  reg  _T_1192_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_472;
  reg  _T_1192_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_473;
  reg  _T_1192_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_474;
  reg  _T_1192_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_475;
  reg  _T_1202_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_476;
  reg  _T_1202_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_477;
  reg  _T_1202_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_478;
  reg  _T_1202_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_479;
  reg  _T_1212_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_480;
  reg  _T_1212_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_481;
  reg  _T_1212_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_482;
  reg  _T_1212_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_483;
  reg  _T_1222_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_484;
  reg  _T_1222_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_485;
  reg  _T_1222_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_486;
  reg  _T_1222_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_487;
  reg  _T_1232_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_488;
  reg  _T_1232_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_489;
  reg  _T_1232_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_490;
  reg  _T_1232_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_491;
  reg  _T_1242_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_492;
  reg  _T_1242_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_493;
  reg  _T_1242_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_494;
  reg  _T_1242_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_495;
  reg  _T_1252_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_496;
  reg  _T_1252_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_497;
  reg  _T_1252_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_498;
  reg  _T_1252_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_499;
  reg  _T_1262_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_500;
  reg  _T_1262_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_501;
  reg  _T_1262_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_502;
  reg  _T_1262_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_503;
  reg  _T_1272_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_504;
  reg  _T_1272_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_505;
  reg  _T_1272_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_506;
  reg  _T_1272_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_507;
  wire  _T_1273 = MultiDimTime_io_index_1 == 18'h16; // @[pearray.scala 182:41]
  wire  _T_1275 = _T_1273 & _T_4; // @[pearray.scala 182:67]
  reg  _T_1282_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_508;
  reg  _T_1282_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_509;
  reg  _T_1282_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_510;
  reg  _T_1282_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_511;
  reg  _T_1292_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_512;
  reg  _T_1292_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_513;
  reg  _T_1292_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_514;
  reg  _T_1292_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_515;
  reg  _T_1302_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_516;
  reg  _T_1302_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_517;
  reg  _T_1302_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_518;
  reg  _T_1302_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_519;
  reg  _T_1312_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_520;
  reg  _T_1312_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_521;
  reg  _T_1312_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_522;
  reg  _T_1312_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_523;
  reg  _T_1322_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_524;
  reg  _T_1322_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_525;
  reg  _T_1322_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_526;
  reg  _T_1322_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_527;
  reg  _T_1332_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_528;
  reg  _T_1332_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_529;
  reg  _T_1332_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_530;
  reg  _T_1332_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_531;
  reg  _T_1342_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_532;
  reg  _T_1342_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_533;
  reg  _T_1342_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_534;
  reg  _T_1342_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_535;
  reg  _T_1352_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_536;
  reg  _T_1352_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_537;
  reg  _T_1352_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_538;
  reg  _T_1352_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_539;
  reg  _T_1362_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_540;
  reg  _T_1362_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_541;
  reg  _T_1362_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_542;
  reg  _T_1362_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_543;
  reg  _T_1372_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_544;
  reg  _T_1372_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_545;
  reg  _T_1372_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_546;
  reg  _T_1372_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_547;
  reg  _T_1382_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_548;
  reg  _T_1382_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_549;
  reg  _T_1382_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_550;
  reg  _T_1382_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_551;
  reg  _T_1392_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_552;
  reg  _T_1392_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_553;
  reg  _T_1392_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_554;
  reg  _T_1392_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_555;
  reg  _T_1402_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_556;
  reg  _T_1402_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_557;
  reg  _T_1402_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_558;
  reg  _T_1402_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_559;
  reg  _T_1412_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_560;
  reg  _T_1412_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_561;
  reg  _T_1412_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_562;
  reg  _T_1412_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_563;
  reg  _T_1422_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_564;
  reg  _T_1422_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_565;
  reg  _T_1422_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_566;
  reg  _T_1422_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_567;
  reg  _T_1432_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_568;
  reg  _T_1432_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_569;
  reg  _T_1432_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_570;
  reg  _T_1432_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_571;
  wire  _T_1433 = MultiDimTime_io_index_1 == 18'h17; // @[pearray.scala 182:41]
  wire  _T_1435 = _T_1433 & _T_4; // @[pearray.scala 182:67]
  reg  _T_1442_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_572;
  reg  _T_1442_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_573;
  reg  _T_1442_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_574;
  reg  _T_1442_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_575;
  reg  _T_1452_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_576;
  reg  _T_1452_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_577;
  reg  _T_1452_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_578;
  reg  _T_1452_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_579;
  reg  _T_1462_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_580;
  reg  _T_1462_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_581;
  reg  _T_1462_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_582;
  reg  _T_1462_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_583;
  reg  _T_1472_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_584;
  reg  _T_1472_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_585;
  reg  _T_1472_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_586;
  reg  _T_1472_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_587;
  reg  _T_1482_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_588;
  reg  _T_1482_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_589;
  reg  _T_1482_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_590;
  reg  _T_1482_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_591;
  reg  _T_1492_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_592;
  reg  _T_1492_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_593;
  reg  _T_1492_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_594;
  reg  _T_1492_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_595;
  reg  _T_1502_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_596;
  reg  _T_1502_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_597;
  reg  _T_1502_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_598;
  reg  _T_1502_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_599;
  reg  _T_1512_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_600;
  reg  _T_1512_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_601;
  reg  _T_1512_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_602;
  reg  _T_1512_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_603;
  reg  _T_1522_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_604;
  reg  _T_1522_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_605;
  reg  _T_1522_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_606;
  reg  _T_1522_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_607;
  reg  _T_1532_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_608;
  reg  _T_1532_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_609;
  reg  _T_1532_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_610;
  reg  _T_1532_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_611;
  reg  _T_1542_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_612;
  reg  _T_1542_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_613;
  reg  _T_1542_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_614;
  reg  _T_1542_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_615;
  reg  _T_1552_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_616;
  reg  _T_1552_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_617;
  reg  _T_1552_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_618;
  reg  _T_1552_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_619;
  reg  _T_1562_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_620;
  reg  _T_1562_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_621;
  reg  _T_1562_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_622;
  reg  _T_1562_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_623;
  reg  _T_1572_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_624;
  reg  _T_1572_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_625;
  reg  _T_1572_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_626;
  reg  _T_1572_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_627;
  reg  _T_1582_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_628;
  reg  _T_1582_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_629;
  reg  _T_1582_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_630;
  reg  _T_1582_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_631;
  reg  _T_1592_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_632;
  reg  _T_1592_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_633;
  reg  _T_1592_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_634;
  reg  _T_1592_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_635;
  wire  _T_1593 = MultiDimTime_io_index_1 == 18'h18; // @[pearray.scala 182:41]
  wire  _T_1595 = _T_1593 & _T_4; // @[pearray.scala 182:67]
  reg  _T_1602_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_636;
  reg  _T_1602_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_637;
  reg  _T_1602_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_638;
  reg  _T_1602_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_639;
  reg  _T_1612_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_640;
  reg  _T_1612_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_641;
  reg  _T_1612_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_642;
  reg  _T_1612_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_643;
  reg  _T_1622_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_644;
  reg  _T_1622_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_645;
  reg  _T_1622_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_646;
  reg  _T_1622_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_647;
  reg  _T_1632_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_648;
  reg  _T_1632_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_649;
  reg  _T_1632_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_650;
  reg  _T_1632_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_651;
  reg  _T_1642_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_652;
  reg  _T_1642_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_653;
  reg  _T_1642_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_654;
  reg  _T_1642_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_655;
  reg  _T_1652_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_656;
  reg  _T_1652_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_657;
  reg  _T_1652_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_658;
  reg  _T_1652_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_659;
  reg  _T_1662_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_660;
  reg  _T_1662_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_661;
  reg  _T_1662_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_662;
  reg  _T_1662_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_663;
  reg  _T_1672_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_664;
  reg  _T_1672_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_665;
  reg  _T_1672_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_666;
  reg  _T_1672_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_667;
  reg  _T_1682_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_668;
  reg  _T_1682_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_669;
  reg  _T_1682_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_670;
  reg  _T_1682_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_671;
  reg  _T_1692_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_672;
  reg  _T_1692_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_673;
  reg  _T_1692_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_674;
  reg  _T_1692_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_675;
  reg  _T_1702_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_676;
  reg  _T_1702_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_677;
  reg  _T_1702_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_678;
  reg  _T_1702_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_679;
  reg  _T_1712_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_680;
  reg  _T_1712_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_681;
  reg  _T_1712_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_682;
  reg  _T_1712_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_683;
  reg  _T_1722_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_684;
  reg  _T_1722_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_685;
  reg  _T_1722_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_686;
  reg  _T_1722_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_687;
  reg  _T_1732_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_688;
  reg  _T_1732_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_689;
  reg  _T_1732_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_690;
  reg  _T_1732_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_691;
  reg  _T_1742_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_692;
  reg  _T_1742_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_693;
  reg  _T_1742_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_694;
  reg  _T_1742_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_695;
  reg  _T_1752_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_696;
  reg  _T_1752_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_697;
  reg  _T_1752_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_698;
  reg  _T_1752_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_699;
  wire  _T_1753 = MultiDimTime_io_index_1 == 18'h19; // @[pearray.scala 182:41]
  wire  _T_1755 = _T_1753 & _T_4; // @[pearray.scala 182:67]
  reg  _T_1762_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_700;
  reg  _T_1762_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_701;
  reg  _T_1762_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_702;
  reg  _T_1762_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_703;
  reg  _T_1772_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_704;
  reg  _T_1772_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_705;
  reg  _T_1772_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_706;
  reg  _T_1772_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_707;
  reg  _T_1782_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_708;
  reg  _T_1782_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_709;
  reg  _T_1782_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_710;
  reg  _T_1782_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_711;
  reg  _T_1792_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_712;
  reg  _T_1792_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_713;
  reg  _T_1792_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_714;
  reg  _T_1792_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_715;
  reg  _T_1802_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_716;
  reg  _T_1802_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_717;
  reg  _T_1802_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_718;
  reg  _T_1802_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_719;
  reg  _T_1812_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_720;
  reg  _T_1812_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_721;
  reg  _T_1812_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_722;
  reg  _T_1812_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_723;
  reg  _T_1822_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_724;
  reg  _T_1822_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_725;
  reg  _T_1822_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_726;
  reg  _T_1822_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_727;
  reg  _T_1832_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_728;
  reg  _T_1832_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_729;
  reg  _T_1832_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_730;
  reg  _T_1832_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_731;
  reg  _T_1842_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_732;
  reg  _T_1842_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_733;
  reg  _T_1842_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_734;
  reg  _T_1842_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_735;
  reg  _T_1852_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_736;
  reg  _T_1852_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_737;
  reg  _T_1852_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_738;
  reg  _T_1852_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_739;
  reg  _T_1862_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_740;
  reg  _T_1862_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_741;
  reg  _T_1862_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_742;
  reg  _T_1862_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_743;
  reg  _T_1872_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_744;
  reg  _T_1872_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_745;
  reg  _T_1872_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_746;
  reg  _T_1872_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_747;
  reg  _T_1882_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_748;
  reg  _T_1882_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_749;
  reg  _T_1882_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_750;
  reg  _T_1882_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_751;
  reg  _T_1892_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_752;
  reg  _T_1892_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_753;
  reg  _T_1892_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_754;
  reg  _T_1892_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_755;
  reg  _T_1902_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_756;
  reg  _T_1902_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_757;
  reg  _T_1902_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_758;
  reg  _T_1902_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_759;
  reg  _T_1912_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_760;
  reg  _T_1912_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_761;
  reg  _T_1912_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_762;
  reg  _T_1912_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_763;
  wire  _T_1913 = MultiDimTime_io_index_1 == 18'h1a; // @[pearray.scala 182:41]
  wire  _T_1915 = _T_1913 & _T_4; // @[pearray.scala 182:67]
  reg  _T_1922_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_764;
  reg  _T_1922_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_765;
  reg  _T_1922_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_766;
  reg  _T_1922_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_767;
  reg  _T_1932_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_768;
  reg  _T_1932_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_769;
  reg  _T_1932_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_770;
  reg  _T_1932_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_771;
  reg  _T_1942_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_772;
  reg  _T_1942_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_773;
  reg  _T_1942_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_774;
  reg  _T_1942_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_775;
  reg  _T_1952_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_776;
  reg  _T_1952_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_777;
  reg  _T_1952_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_778;
  reg  _T_1952_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_779;
  reg  _T_1962_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_780;
  reg  _T_1962_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_781;
  reg  _T_1962_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_782;
  reg  _T_1962_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_783;
  reg  _T_1972_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_784;
  reg  _T_1972_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_785;
  reg  _T_1972_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_786;
  reg  _T_1972_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_787;
  reg  _T_1982_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_788;
  reg  _T_1982_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_789;
  reg  _T_1982_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_790;
  reg  _T_1982_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_791;
  reg  _T_1992_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_792;
  reg  _T_1992_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_793;
  reg  _T_1992_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_794;
  reg  _T_1992_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_795;
  reg  _T_2002_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_796;
  reg  _T_2002_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_797;
  reg  _T_2002_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_798;
  reg  _T_2002_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_799;
  reg  _T_2012_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_800;
  reg  _T_2012_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_801;
  reg  _T_2012_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_802;
  reg  _T_2012_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_803;
  reg  _T_2022_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_804;
  reg  _T_2022_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_805;
  reg  _T_2022_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_806;
  reg  _T_2022_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_807;
  reg  _T_2032_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_808;
  reg  _T_2032_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_809;
  reg  _T_2032_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_810;
  reg  _T_2032_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_811;
  reg  _T_2042_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_812;
  reg  _T_2042_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_813;
  reg  _T_2042_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_814;
  reg  _T_2042_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_815;
  reg  _T_2052_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_816;
  reg  _T_2052_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_817;
  reg  _T_2052_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_818;
  reg  _T_2052_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_819;
  reg  _T_2062_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_820;
  reg  _T_2062_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_821;
  reg  _T_2062_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_822;
  reg  _T_2062_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_823;
  reg  _T_2072_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_824;
  reg  _T_2072_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_825;
  reg  _T_2072_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_826;
  reg  _T_2072_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_827;
  wire  _T_2073 = MultiDimTime_io_index_1 == 18'h1b; // @[pearray.scala 182:41]
  wire  _T_2075 = _T_2073 & _T_4; // @[pearray.scala 182:67]
  reg  _T_2082_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_828;
  reg  _T_2082_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_829;
  reg  _T_2082_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_830;
  reg  _T_2082_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_831;
  reg  _T_2092_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_832;
  reg  _T_2092_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_833;
  reg  _T_2092_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_834;
  reg  _T_2092_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_835;
  reg  _T_2102_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_836;
  reg  _T_2102_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_837;
  reg  _T_2102_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_838;
  reg  _T_2102_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_839;
  reg  _T_2112_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_840;
  reg  _T_2112_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_841;
  reg  _T_2112_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_842;
  reg  _T_2112_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_843;
  reg  _T_2122_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_844;
  reg  _T_2122_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_845;
  reg  _T_2122_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_846;
  reg  _T_2122_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_847;
  reg  _T_2132_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_848;
  reg  _T_2132_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_849;
  reg  _T_2132_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_850;
  reg  _T_2132_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_851;
  reg  _T_2142_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_852;
  reg  _T_2142_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_853;
  reg  _T_2142_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_854;
  reg  _T_2142_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_855;
  reg  _T_2152_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_856;
  reg  _T_2152_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_857;
  reg  _T_2152_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_858;
  reg  _T_2152_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_859;
  reg  _T_2162_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_860;
  reg  _T_2162_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_861;
  reg  _T_2162_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_862;
  reg  _T_2162_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_863;
  reg  _T_2172_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_864;
  reg  _T_2172_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_865;
  reg  _T_2172_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_866;
  reg  _T_2172_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_867;
  reg  _T_2182_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_868;
  reg  _T_2182_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_869;
  reg  _T_2182_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_870;
  reg  _T_2182_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_871;
  reg  _T_2192_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_872;
  reg  _T_2192_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_873;
  reg  _T_2192_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_874;
  reg  _T_2192_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_875;
  reg  _T_2202_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_876;
  reg  _T_2202_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_877;
  reg  _T_2202_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_878;
  reg  _T_2202_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_879;
  reg  _T_2212_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_880;
  reg  _T_2212_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_881;
  reg  _T_2212_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_882;
  reg  _T_2212_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_883;
  reg  _T_2222_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_884;
  reg  _T_2222_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_885;
  reg  _T_2222_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_886;
  reg  _T_2222_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_887;
  reg  _T_2232_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_888;
  reg  _T_2232_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_889;
  reg  _T_2232_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_890;
  reg  _T_2232_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_891;
  wire  _T_2233 = MultiDimTime_io_index_1 == 18'h1c; // @[pearray.scala 182:41]
  wire  _T_2235 = _T_2233 & _T_4; // @[pearray.scala 182:67]
  reg  _T_2242_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_892;
  reg  _T_2242_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_893;
  reg  _T_2242_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_894;
  reg  _T_2242_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_895;
  reg  _T_2252_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_896;
  reg  _T_2252_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_897;
  reg  _T_2252_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_898;
  reg  _T_2252_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_899;
  reg  _T_2262_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_900;
  reg  _T_2262_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_901;
  reg  _T_2262_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_902;
  reg  _T_2262_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_903;
  reg  _T_2272_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_904;
  reg  _T_2272_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_905;
  reg  _T_2272_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_906;
  reg  _T_2272_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_907;
  reg  _T_2282_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_908;
  reg  _T_2282_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_909;
  reg  _T_2282_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_910;
  reg  _T_2282_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_911;
  reg  _T_2292_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_912;
  reg  _T_2292_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_913;
  reg  _T_2292_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_914;
  reg  _T_2292_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_915;
  reg  _T_2302_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_916;
  reg  _T_2302_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_917;
  reg  _T_2302_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_918;
  reg  _T_2302_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_919;
  reg  _T_2312_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_920;
  reg  _T_2312_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_921;
  reg  _T_2312_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_922;
  reg  _T_2312_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_923;
  reg  _T_2322_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_924;
  reg  _T_2322_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_925;
  reg  _T_2322_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_926;
  reg  _T_2322_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_927;
  reg  _T_2332_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_928;
  reg  _T_2332_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_929;
  reg  _T_2332_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_930;
  reg  _T_2332_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_931;
  reg  _T_2342_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_932;
  reg  _T_2342_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_933;
  reg  _T_2342_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_934;
  reg  _T_2342_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_935;
  reg  _T_2352_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_936;
  reg  _T_2352_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_937;
  reg  _T_2352_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_938;
  reg  _T_2352_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_939;
  reg  _T_2362_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_940;
  reg  _T_2362_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_941;
  reg  _T_2362_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_942;
  reg  _T_2362_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_943;
  reg  _T_2372_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_944;
  reg  _T_2372_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_945;
  reg  _T_2372_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_946;
  reg  _T_2372_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_947;
  reg  _T_2382_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_948;
  reg  _T_2382_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_949;
  reg  _T_2382_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_950;
  reg  _T_2382_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_951;
  reg  _T_2392_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_952;
  reg  _T_2392_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_953;
  reg  _T_2392_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_954;
  reg  _T_2392_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_955;
  wire  _T_2393 = MultiDimTime_io_index_1 == 18'h1d; // @[pearray.scala 182:41]
  wire  _T_2395 = _T_2393 & _T_4; // @[pearray.scala 182:67]
  reg  _T_2402_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_956;
  reg  _T_2402_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_957;
  reg  _T_2402_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_958;
  reg  _T_2402_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_959;
  reg  _T_2412_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_960;
  reg  _T_2412_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_961;
  reg  _T_2412_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_962;
  reg  _T_2412_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_963;
  reg  _T_2422_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_964;
  reg  _T_2422_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_965;
  reg  _T_2422_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_966;
  reg  _T_2422_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_967;
  reg  _T_2432_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_968;
  reg  _T_2432_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_969;
  reg  _T_2432_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_970;
  reg  _T_2432_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_971;
  reg  _T_2442_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_972;
  reg  _T_2442_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_973;
  reg  _T_2442_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_974;
  reg  _T_2442_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_975;
  reg  _T_2452_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_976;
  reg  _T_2452_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_977;
  reg  _T_2452_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_978;
  reg  _T_2452_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_979;
  reg  _T_2462_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_980;
  reg  _T_2462_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_981;
  reg  _T_2462_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_982;
  reg  _T_2462_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_983;
  reg  _T_2472_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_984;
  reg  _T_2472_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_985;
  reg  _T_2472_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_986;
  reg  _T_2472_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_987;
  reg  _T_2482_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_988;
  reg  _T_2482_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_989;
  reg  _T_2482_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_990;
  reg  _T_2482_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_991;
  reg  _T_2492_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_992;
  reg  _T_2492_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_993;
  reg  _T_2492_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_994;
  reg  _T_2492_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_995;
  reg  _T_2502_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_996;
  reg  _T_2502_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_997;
  reg  _T_2502_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_998;
  reg  _T_2502_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_999;
  reg  _T_2512_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1000;
  reg  _T_2512_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1001;
  reg  _T_2512_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1002;
  reg  _T_2512_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1003;
  reg  _T_2522_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1004;
  reg  _T_2522_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1005;
  reg  _T_2522_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1006;
  reg  _T_2522_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1007;
  reg  _T_2532_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1008;
  reg  _T_2532_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1009;
  reg  _T_2532_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1010;
  reg  _T_2532_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1011;
  reg  _T_2542_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1012;
  reg  _T_2542_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1013;
  reg  _T_2542_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1014;
  reg  _T_2542_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1015;
  reg  _T_2552_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1016;
  reg  _T_2552_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1017;
  reg  _T_2552_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1018;
  reg  _T_2552_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1019;
  wire  _T_2553 = MultiDimTime_io_index_1 == 18'h1e; // @[pearray.scala 182:41]
  wire  _T_2555 = _T_2553 & _T_4; // @[pearray.scala 182:67]
  reg  _T_2562_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1020;
  reg  _T_2562_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1021;
  reg  _T_2562_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1022;
  reg  _T_2562_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1023;
  wire  _T_2569 = MultiDimTime_io_index_1 < 18'h10; // @[pearray.scala 252:134]
  wire  _T_2570 = io_exec_valid & _T_2569; // @[pearray.scala 252:112]
  reg  _T_2575_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1024;
  reg  _T_2575_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1025;
  reg  _T_2575_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1026;
  wire  _T_2576 = MultiDimTime_io_index_1 >= 18'h1; // @[pearray.scala 252:82]
  wire  _T_2577 = io_exec_valid & _T_2576; // @[pearray.scala 252:60]
  wire  _T_2578 = MultiDimTime_io_index_1 < 18'h11; // @[pearray.scala 252:134]
  wire  _T_2579 = _T_2577 & _T_2578; // @[pearray.scala 252:112]
  reg  _T_2584_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1027;
  reg  _T_2584_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1028;
  reg  _T_2584_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1029;
  wire  _T_2585 = MultiDimTime_io_index_1 >= 18'h2; // @[pearray.scala 252:82]
  wire  _T_2586 = io_exec_valid & _T_2585; // @[pearray.scala 252:60]
  wire  _T_2587 = MultiDimTime_io_index_1 < 18'h12; // @[pearray.scala 252:134]
  wire  _T_2588 = _T_2586 & _T_2587; // @[pearray.scala 252:112]
  reg  _T_2593_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1030;
  reg  _T_2593_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1031;
  reg  _T_2593_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1032;
  wire  _T_2594 = MultiDimTime_io_index_1 >= 18'h3; // @[pearray.scala 252:82]
  wire  _T_2595 = io_exec_valid & _T_2594; // @[pearray.scala 252:60]
  wire  _T_2596 = MultiDimTime_io_index_1 < 18'h13; // @[pearray.scala 252:134]
  wire  _T_2597 = _T_2595 & _T_2596; // @[pearray.scala 252:112]
  reg  _T_2602_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1033;
  reg  _T_2602_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1034;
  reg  _T_2602_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1035;
  wire  _T_2603 = MultiDimTime_io_index_1 >= 18'h4; // @[pearray.scala 252:82]
  wire  _T_2604 = io_exec_valid & _T_2603; // @[pearray.scala 252:60]
  wire  _T_2605 = MultiDimTime_io_index_1 < 18'h14; // @[pearray.scala 252:134]
  wire  _T_2606 = _T_2604 & _T_2605; // @[pearray.scala 252:112]
  reg  _T_2611_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1036;
  reg  _T_2611_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1037;
  reg  _T_2611_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1038;
  wire  _T_2612 = MultiDimTime_io_index_1 >= 18'h5; // @[pearray.scala 252:82]
  wire  _T_2613 = io_exec_valid & _T_2612; // @[pearray.scala 252:60]
  wire  _T_2614 = MultiDimTime_io_index_1 < 18'h15; // @[pearray.scala 252:134]
  wire  _T_2615 = _T_2613 & _T_2614; // @[pearray.scala 252:112]
  reg  _T_2620_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1039;
  reg  _T_2620_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1040;
  reg  _T_2620_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1041;
  wire  _T_2621 = MultiDimTime_io_index_1 >= 18'h6; // @[pearray.scala 252:82]
  wire  _T_2622 = io_exec_valid & _T_2621; // @[pearray.scala 252:60]
  wire  _T_2623 = MultiDimTime_io_index_1 < 18'h16; // @[pearray.scala 252:134]
  wire  _T_2624 = _T_2622 & _T_2623; // @[pearray.scala 252:112]
  reg  _T_2629_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1042;
  reg  _T_2629_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1043;
  reg  _T_2629_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1044;
  wire  _T_2630 = MultiDimTime_io_index_1 >= 18'h7; // @[pearray.scala 252:82]
  wire  _T_2631 = io_exec_valid & _T_2630; // @[pearray.scala 252:60]
  wire  _T_2632 = MultiDimTime_io_index_1 < 18'h17; // @[pearray.scala 252:134]
  wire  _T_2633 = _T_2631 & _T_2632; // @[pearray.scala 252:112]
  reg  _T_2638_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1045;
  reg  _T_2638_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1046;
  reg  _T_2638_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1047;
  wire  _T_2639 = MultiDimTime_io_index_1 >= 18'h8; // @[pearray.scala 252:82]
  wire  _T_2640 = io_exec_valid & _T_2639; // @[pearray.scala 252:60]
  wire  _T_2641 = MultiDimTime_io_index_1 < 18'h18; // @[pearray.scala 252:134]
  wire  _T_2642 = _T_2640 & _T_2641; // @[pearray.scala 252:112]
  reg  _T_2647_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1048;
  reg  _T_2647_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1049;
  reg  _T_2647_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1050;
  wire  _T_2648 = MultiDimTime_io_index_1 >= 18'h9; // @[pearray.scala 252:82]
  wire  _T_2649 = io_exec_valid & _T_2648; // @[pearray.scala 252:60]
  wire  _T_2650 = MultiDimTime_io_index_1 < 18'h19; // @[pearray.scala 252:134]
  wire  _T_2651 = _T_2649 & _T_2650; // @[pearray.scala 252:112]
  reg  _T_2656_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1051;
  reg  _T_2656_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1052;
  reg  _T_2656_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1053;
  wire  _T_2657 = MultiDimTime_io_index_1 >= 18'ha; // @[pearray.scala 252:82]
  wire  _T_2658 = io_exec_valid & _T_2657; // @[pearray.scala 252:60]
  wire  _T_2659 = MultiDimTime_io_index_1 < 18'h1a; // @[pearray.scala 252:134]
  wire  _T_2660 = _T_2658 & _T_2659; // @[pearray.scala 252:112]
  reg  _T_2665_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1054;
  reg  _T_2665_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1055;
  reg  _T_2665_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1056;
  wire  _T_2666 = MultiDimTime_io_index_1 >= 18'hb; // @[pearray.scala 252:82]
  wire  _T_2667 = io_exec_valid & _T_2666; // @[pearray.scala 252:60]
  wire  _T_2668 = MultiDimTime_io_index_1 < 18'h1b; // @[pearray.scala 252:134]
  wire  _T_2669 = _T_2667 & _T_2668; // @[pearray.scala 252:112]
  reg  _T_2674_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1057;
  reg  _T_2674_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1058;
  reg  _T_2674_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1059;
  wire  _T_2675 = MultiDimTime_io_index_1 >= 18'hc; // @[pearray.scala 252:82]
  wire  _T_2676 = io_exec_valid & _T_2675; // @[pearray.scala 252:60]
  wire  _T_2677 = MultiDimTime_io_index_1 < 18'h1c; // @[pearray.scala 252:134]
  wire  _T_2678 = _T_2676 & _T_2677; // @[pearray.scala 252:112]
  reg  _T_2683_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1060;
  reg  _T_2683_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1061;
  reg  _T_2683_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1062;
  wire  _T_2684 = MultiDimTime_io_index_1 >= 18'hd; // @[pearray.scala 252:82]
  wire  _T_2685 = io_exec_valid & _T_2684; // @[pearray.scala 252:60]
  wire  _T_2686 = MultiDimTime_io_index_1 < 18'h1d; // @[pearray.scala 252:134]
  wire  _T_2687 = _T_2685 & _T_2686; // @[pearray.scala 252:112]
  reg  _T_2692_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1063;
  reg  _T_2692_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1064;
  reg  _T_2692_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1065;
  wire  _T_2693 = MultiDimTime_io_index_1 >= 18'he; // @[pearray.scala 252:82]
  wire  _T_2694 = io_exec_valid & _T_2693; // @[pearray.scala 252:60]
  wire  _T_2695 = MultiDimTime_io_index_1 < 18'h1e; // @[pearray.scala 252:134]
  wire  _T_2696 = _T_2694 & _T_2695; // @[pearray.scala 252:112]
  reg  _T_2701_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1066;
  reg  _T_2701_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1067;
  reg  _T_2701_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1068;
  wire  _T_2702 = MultiDimTime_io_index_1 >= 18'hf; // @[pearray.scala 252:82]
  wire  _T_2703 = io_exec_valid & _T_2702; // @[pearray.scala 252:60]
  wire  _T_2704 = MultiDimTime_io_index_1 < 18'h1f; // @[pearray.scala 252:134]
  wire  _T_2705 = _T_2703 & _T_2704; // @[pearray.scala 252:112]
  reg  _T_2710_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1069;
  reg  _T_2710_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1070;
  reg  _T_2710_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1071;
  reg  _T_2712_0; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1072;
  reg  _T_2712_1; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1073;
  reg  _T_2712_2; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1074;
  reg  _T_2712_3; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1075;
  reg  _T_2712_4; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1076;
  reg  _T_2712_5; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1077;
  reg  _T_2712_6; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1078;
  reg  _T_2712_7; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1079;
  reg  _T_2712_8; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1080;
  reg  _T_2712_9; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1081;
  reg  _T_2712_10; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1082;
  reg  _T_2712_11; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1083;
  reg  _T_2712_12; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1084;
  reg  _T_2712_13; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1085;
  reg  _T_2712_14; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1086;
  reg  _T_2712_15; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1087;
  reg  _T_2712_16; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1088;
  reg  _T_2712_17; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1089;
  reg  _T_2712_18; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1090;
  reg  _T_2712_19; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1091;
  reg  _T_2712_20; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1092;
  reg  _T_2712_21; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1093;
  reg  _T_2712_22; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1094;
  reg  _T_2712_23; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1095;
  reg  _T_2712_24; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1096;
  reg  _T_2712_25; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1097;
  reg  _T_2712_26; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1098;
  reg  _T_2712_27; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1099;
  reg  _T_2712_28; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1100;
  reg  _T_2712_29; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1101;
  reg  _T_2712_30; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1102;
  reg  _T_2712_31; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1103;
  reg  _T_2712_32; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1104;
  reg  _T_2712_33; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1105;
  reg  _T_2712_34; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1106;
  reg  _T_2712_35; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1107;
  reg  _T_2712_36; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1108;
  reg  _T_2712_37; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1109;
  reg  _T_2712_38; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1110;
  reg  _T_2712_39; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1111;
  reg  _T_2712_40; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1112;
  reg  _T_2712_41; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1113;
  reg  _T_2712_42; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1114;
  reg  _T_2712_43; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1115;
  reg  _T_2712_44; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1116;
  reg  _T_2712_45; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1117;
  reg  _T_2712_46; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1118;
  reg  _T_2712_47; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1119;
  reg  _T_2712_48; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1120;
  reg  _T_2712_49; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1121;
  reg  _T_2712_50; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1122;
  reg  _T_2712_51; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1123;
  reg  _T_2712_52; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1124;
  reg  _T_2712_53; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1125;
  reg  _T_2712_54; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1126;
  reg  _T_2712_55; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1127;
  reg  _T_2712_56; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1128;
  reg  _T_2712_57; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1129;
  reg  _T_2712_58; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1130;
  reg  _T_2712_59; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1131;
  reg  _T_2712_60; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1132;
  reg  _T_2712_61; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1133;
  reg  _T_2712_62; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1134;
  reg  _T_2712_63; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1135;
  reg  _T_2712_64; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1136;
  reg  _T_2712_65; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1137;
  reg  _T_2712_66; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1138;
  reg  _T_2712_67; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1139;
  reg  _T_2712_68; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1140;
  reg  _T_2712_69; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1141;
  reg  _T_2712_70; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1142;
  reg  _T_2712_71; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1143;
  reg  _T_2712_72; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1144;
  reg  _T_2712_73; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1145;
  reg  _T_2712_74; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1146;
  reg  _T_2712_75; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1147;
  reg  _T_2712_76; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1148;
  reg  _T_2712_77; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1149;
  reg  _T_2712_78; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1150;
  reg  _T_2712_79; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1151;
  reg  _T_2712_80; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1152;
  reg  _T_2712_81; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1153;
  reg  _T_2712_82; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1154;
  reg  _T_2712_83; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1155;
  reg  _T_2712_84; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1156;
  reg  _T_2712_85; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1157;
  reg  _T_2712_86; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1158;
  reg  _T_2712_87; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1159;
  reg  _T_2712_88; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1160;
  reg  _T_2712_89; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1161;
  reg  _T_2712_90; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1162;
  reg  _T_2712_91; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1163;
  reg  _T_2712_92; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1164;
  reg  _T_2712_93; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1165;
  reg  _T_2712_94; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1166;
  reg  _T_2712_95; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1167;
  reg  _T_2712_96; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1168;
  reg  _T_2712_97; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1169;
  reg  _T_2712_98; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1170;
  reg  _T_2712_99; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1171;
  reg  _T_2712_100; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1172;
  reg  _T_2712_101; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1173;
  reg  _T_2712_102; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1174;
  reg  _T_2712_103; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1175;
  reg  _T_2712_104; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1176;
  reg  _T_2712_105; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1177;
  reg  _T_2712_106; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1178;
  reg  _T_2712_107; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1179;
  reg  _T_2712_108; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1180;
  reg  _T_2712_109; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1181;
  reg  _T_2712_110; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1182;
  reg  _T_2712_111; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1183;
  reg  _T_2712_112; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1184;
  reg  _T_2712_113; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1185;
  reg  _T_2712_114; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1186;
  reg  _T_2712_115; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1187;
  reg  _T_2712_116; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1188;
  reg  _T_2712_117; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1189;
  reg  _T_2712_118; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1190;
  reg  _T_2712_119; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1191;
  reg  _T_2712_120; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1192;
  reg  _T_2712_121; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1193;
  reg  _T_2712_122; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1194;
  reg  _T_2712_123; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1195;
  reg  _T_2712_124; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1196;
  reg  _T_2712_125; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1197;
  reg  _T_2712_126; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1198;
  reg  _T_2712_127; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1199;
  reg  _T_2712_128; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1200;
  reg  _T_2712_129; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1201;
  reg  _T_2712_130; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1202;
  reg  _T_2712_131; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1203;
  reg  _T_2712_132; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1204;
  reg  _T_2712_133; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1205;
  reg  _T_2712_134; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1206;
  reg  _T_2712_135; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1207;
  reg  _T_2712_136; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1208;
  reg  _T_2712_137; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1209;
  reg  _T_2712_138; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1210;
  reg  _T_2712_139; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1211;
  reg  _T_2712_140; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1212;
  reg  _T_2712_141; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1213;
  reg  _T_2712_142; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1214;
  reg  _T_2712_143; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1215;
  reg  _T_2712_144; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1216;
  reg  _T_2712_145; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1217;
  reg  _T_2712_146; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1218;
  reg  _T_2712_147; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1219;
  reg  _T_2712_148; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1220;
  reg  _T_2712_149; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1221;
  reg  _T_2712_150; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1222;
  reg  _T_2712_151; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1223;
  reg  _T_2712_152; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1224;
  reg  _T_2712_153; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1225;
  reg  _T_2712_154; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1226;
  reg  _T_2712_155; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1227;
  reg  _T_2712_156; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1228;
  reg  _T_2712_157; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1229;
  reg  _T_2712_158; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1230;
  reg  _T_2712_159; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1231;
  reg  _T_2712_160; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1232;
  reg  _T_2712_161; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1233;
  reg  _T_2712_162; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1234;
  reg  _T_2712_163; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1235;
  reg  _T_2712_164; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1236;
  reg  _T_2712_165; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1237;
  reg  _T_2712_166; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1238;
  reg  _T_2712_167; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1239;
  reg  _T_2712_168; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1240;
  reg  _T_2712_169; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1241;
  reg  _T_2712_170; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1242;
  reg  _T_2712_171; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1243;
  reg  _T_2712_172; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1244;
  reg  _T_2712_173; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1245;
  reg  _T_2712_174; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1246;
  reg  _T_2712_175; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1247;
  reg  _T_2712_176; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1248;
  reg  _T_2712_177; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1249;
  reg  _T_2712_178; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1250;
  reg  _T_2712_179; // @[pearray.scala 225:27]
  reg [31:0] _RAND_1251;
  MultiDimTime MultiDimTime ( // @[pearray.scala 63:25]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_out_3(MultiDimTime_io_out_3),
    .io_out_4(MultiDimTime_io_out_4),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2),
    .io_index_3(MultiDimTime_io_index_3)
  );
  PE PE ( // @[pearray.scala 103:13]
    .clock(PE_clock),
    .reset(PE_reset),
    .io_data_2_in_valid(PE_io_data_2_in_valid),
    .io_data_2_in_bits(PE_io_data_2_in_bits),
    .io_data_2_out_valid(PE_io_data_2_out_valid),
    .io_data_2_out_bits(PE_io_data_2_out_bits),
    .io_data_1_in_valid(PE_io_data_1_in_valid),
    .io_data_1_in_bits(PE_io_data_1_in_bits),
    .io_data_1_out_valid(PE_io_data_1_out_valid),
    .io_data_1_out_bits(PE_io_data_1_out_bits),
    .io_data_0_in_valid(PE_io_data_0_in_valid),
    .io_data_0_in_bits(PE_io_data_0_in_bits),
    .io_data_0_out_valid(PE_io_data_0_out_valid),
    .io_data_0_out_bits(PE_io_data_0_out_bits),
    .io_sig_stat2trans(PE_io_sig_stat2trans)
  );
  PE PE_1 ( // @[pearray.scala 103:13]
    .clock(PE_1_clock),
    .reset(PE_1_reset),
    .io_data_2_in_valid(PE_1_io_data_2_in_valid),
    .io_data_2_in_bits(PE_1_io_data_2_in_bits),
    .io_data_2_out_valid(PE_1_io_data_2_out_valid),
    .io_data_2_out_bits(PE_1_io_data_2_out_bits),
    .io_data_1_in_valid(PE_1_io_data_1_in_valid),
    .io_data_1_in_bits(PE_1_io_data_1_in_bits),
    .io_data_1_out_valid(PE_1_io_data_1_out_valid),
    .io_data_1_out_bits(PE_1_io_data_1_out_bits),
    .io_data_0_in_valid(PE_1_io_data_0_in_valid),
    .io_data_0_in_bits(PE_1_io_data_0_in_bits),
    .io_data_0_out_valid(PE_1_io_data_0_out_valid),
    .io_data_0_out_bits(PE_1_io_data_0_out_bits),
    .io_sig_stat2trans(PE_1_io_sig_stat2trans)
  );
  PE PE_2 ( // @[pearray.scala 103:13]
    .clock(PE_2_clock),
    .reset(PE_2_reset),
    .io_data_2_in_valid(PE_2_io_data_2_in_valid),
    .io_data_2_in_bits(PE_2_io_data_2_in_bits),
    .io_data_2_out_valid(PE_2_io_data_2_out_valid),
    .io_data_2_out_bits(PE_2_io_data_2_out_bits),
    .io_data_1_in_valid(PE_2_io_data_1_in_valid),
    .io_data_1_in_bits(PE_2_io_data_1_in_bits),
    .io_data_1_out_valid(PE_2_io_data_1_out_valid),
    .io_data_1_out_bits(PE_2_io_data_1_out_bits),
    .io_data_0_in_valid(PE_2_io_data_0_in_valid),
    .io_data_0_in_bits(PE_2_io_data_0_in_bits),
    .io_data_0_out_valid(PE_2_io_data_0_out_valid),
    .io_data_0_out_bits(PE_2_io_data_0_out_bits),
    .io_sig_stat2trans(PE_2_io_sig_stat2trans)
  );
  PE PE_3 ( // @[pearray.scala 103:13]
    .clock(PE_3_clock),
    .reset(PE_3_reset),
    .io_data_2_in_valid(PE_3_io_data_2_in_valid),
    .io_data_2_in_bits(PE_3_io_data_2_in_bits),
    .io_data_2_out_valid(PE_3_io_data_2_out_valid),
    .io_data_2_out_bits(PE_3_io_data_2_out_bits),
    .io_data_1_in_valid(PE_3_io_data_1_in_valid),
    .io_data_1_in_bits(PE_3_io_data_1_in_bits),
    .io_data_1_out_valid(PE_3_io_data_1_out_valid),
    .io_data_1_out_bits(PE_3_io_data_1_out_bits),
    .io_data_0_in_valid(PE_3_io_data_0_in_valid),
    .io_data_0_in_bits(PE_3_io_data_0_in_bits),
    .io_data_0_out_valid(PE_3_io_data_0_out_valid),
    .io_data_0_out_bits(PE_3_io_data_0_out_bits),
    .io_sig_stat2trans(PE_3_io_sig_stat2trans)
  );
  PE PE_4 ( // @[pearray.scala 103:13]
    .clock(PE_4_clock),
    .reset(PE_4_reset),
    .io_data_2_in_valid(PE_4_io_data_2_in_valid),
    .io_data_2_in_bits(PE_4_io_data_2_in_bits),
    .io_data_2_out_valid(PE_4_io_data_2_out_valid),
    .io_data_2_out_bits(PE_4_io_data_2_out_bits),
    .io_data_1_in_valid(PE_4_io_data_1_in_valid),
    .io_data_1_in_bits(PE_4_io_data_1_in_bits),
    .io_data_1_out_valid(PE_4_io_data_1_out_valid),
    .io_data_1_out_bits(PE_4_io_data_1_out_bits),
    .io_data_0_in_valid(PE_4_io_data_0_in_valid),
    .io_data_0_in_bits(PE_4_io_data_0_in_bits),
    .io_data_0_out_valid(PE_4_io_data_0_out_valid),
    .io_data_0_out_bits(PE_4_io_data_0_out_bits),
    .io_sig_stat2trans(PE_4_io_sig_stat2trans)
  );
  PE PE_5 ( // @[pearray.scala 103:13]
    .clock(PE_5_clock),
    .reset(PE_5_reset),
    .io_data_2_in_valid(PE_5_io_data_2_in_valid),
    .io_data_2_in_bits(PE_5_io_data_2_in_bits),
    .io_data_2_out_valid(PE_5_io_data_2_out_valid),
    .io_data_2_out_bits(PE_5_io_data_2_out_bits),
    .io_data_1_in_valid(PE_5_io_data_1_in_valid),
    .io_data_1_in_bits(PE_5_io_data_1_in_bits),
    .io_data_1_out_valid(PE_5_io_data_1_out_valid),
    .io_data_1_out_bits(PE_5_io_data_1_out_bits),
    .io_data_0_in_valid(PE_5_io_data_0_in_valid),
    .io_data_0_in_bits(PE_5_io_data_0_in_bits),
    .io_data_0_out_valid(PE_5_io_data_0_out_valid),
    .io_data_0_out_bits(PE_5_io_data_0_out_bits),
    .io_sig_stat2trans(PE_5_io_sig_stat2trans)
  );
  PE PE_6 ( // @[pearray.scala 103:13]
    .clock(PE_6_clock),
    .reset(PE_6_reset),
    .io_data_2_in_valid(PE_6_io_data_2_in_valid),
    .io_data_2_in_bits(PE_6_io_data_2_in_bits),
    .io_data_2_out_valid(PE_6_io_data_2_out_valid),
    .io_data_2_out_bits(PE_6_io_data_2_out_bits),
    .io_data_1_in_valid(PE_6_io_data_1_in_valid),
    .io_data_1_in_bits(PE_6_io_data_1_in_bits),
    .io_data_1_out_valid(PE_6_io_data_1_out_valid),
    .io_data_1_out_bits(PE_6_io_data_1_out_bits),
    .io_data_0_in_valid(PE_6_io_data_0_in_valid),
    .io_data_0_in_bits(PE_6_io_data_0_in_bits),
    .io_data_0_out_valid(PE_6_io_data_0_out_valid),
    .io_data_0_out_bits(PE_6_io_data_0_out_bits),
    .io_sig_stat2trans(PE_6_io_sig_stat2trans)
  );
  PE PE_7 ( // @[pearray.scala 103:13]
    .clock(PE_7_clock),
    .reset(PE_7_reset),
    .io_data_2_in_valid(PE_7_io_data_2_in_valid),
    .io_data_2_in_bits(PE_7_io_data_2_in_bits),
    .io_data_2_out_valid(PE_7_io_data_2_out_valid),
    .io_data_2_out_bits(PE_7_io_data_2_out_bits),
    .io_data_1_in_valid(PE_7_io_data_1_in_valid),
    .io_data_1_in_bits(PE_7_io_data_1_in_bits),
    .io_data_1_out_valid(PE_7_io_data_1_out_valid),
    .io_data_1_out_bits(PE_7_io_data_1_out_bits),
    .io_data_0_in_valid(PE_7_io_data_0_in_valid),
    .io_data_0_in_bits(PE_7_io_data_0_in_bits),
    .io_data_0_out_valid(PE_7_io_data_0_out_valid),
    .io_data_0_out_bits(PE_7_io_data_0_out_bits),
    .io_sig_stat2trans(PE_7_io_sig_stat2trans)
  );
  PE PE_8 ( // @[pearray.scala 103:13]
    .clock(PE_8_clock),
    .reset(PE_8_reset),
    .io_data_2_in_valid(PE_8_io_data_2_in_valid),
    .io_data_2_in_bits(PE_8_io_data_2_in_bits),
    .io_data_2_out_valid(PE_8_io_data_2_out_valid),
    .io_data_2_out_bits(PE_8_io_data_2_out_bits),
    .io_data_1_in_valid(PE_8_io_data_1_in_valid),
    .io_data_1_in_bits(PE_8_io_data_1_in_bits),
    .io_data_1_out_valid(PE_8_io_data_1_out_valid),
    .io_data_1_out_bits(PE_8_io_data_1_out_bits),
    .io_data_0_in_valid(PE_8_io_data_0_in_valid),
    .io_data_0_in_bits(PE_8_io_data_0_in_bits),
    .io_data_0_out_valid(PE_8_io_data_0_out_valid),
    .io_data_0_out_bits(PE_8_io_data_0_out_bits),
    .io_sig_stat2trans(PE_8_io_sig_stat2trans)
  );
  PE PE_9 ( // @[pearray.scala 103:13]
    .clock(PE_9_clock),
    .reset(PE_9_reset),
    .io_data_2_in_valid(PE_9_io_data_2_in_valid),
    .io_data_2_in_bits(PE_9_io_data_2_in_bits),
    .io_data_2_out_valid(PE_9_io_data_2_out_valid),
    .io_data_2_out_bits(PE_9_io_data_2_out_bits),
    .io_data_1_in_valid(PE_9_io_data_1_in_valid),
    .io_data_1_in_bits(PE_9_io_data_1_in_bits),
    .io_data_1_out_valid(PE_9_io_data_1_out_valid),
    .io_data_1_out_bits(PE_9_io_data_1_out_bits),
    .io_data_0_in_valid(PE_9_io_data_0_in_valid),
    .io_data_0_in_bits(PE_9_io_data_0_in_bits),
    .io_data_0_out_valid(PE_9_io_data_0_out_valid),
    .io_data_0_out_bits(PE_9_io_data_0_out_bits),
    .io_sig_stat2trans(PE_9_io_sig_stat2trans)
  );
  PE PE_10 ( // @[pearray.scala 103:13]
    .clock(PE_10_clock),
    .reset(PE_10_reset),
    .io_data_2_in_valid(PE_10_io_data_2_in_valid),
    .io_data_2_in_bits(PE_10_io_data_2_in_bits),
    .io_data_2_out_valid(PE_10_io_data_2_out_valid),
    .io_data_2_out_bits(PE_10_io_data_2_out_bits),
    .io_data_1_in_valid(PE_10_io_data_1_in_valid),
    .io_data_1_in_bits(PE_10_io_data_1_in_bits),
    .io_data_1_out_valid(PE_10_io_data_1_out_valid),
    .io_data_1_out_bits(PE_10_io_data_1_out_bits),
    .io_data_0_in_valid(PE_10_io_data_0_in_valid),
    .io_data_0_in_bits(PE_10_io_data_0_in_bits),
    .io_data_0_out_valid(PE_10_io_data_0_out_valid),
    .io_data_0_out_bits(PE_10_io_data_0_out_bits),
    .io_sig_stat2trans(PE_10_io_sig_stat2trans)
  );
  PE PE_11 ( // @[pearray.scala 103:13]
    .clock(PE_11_clock),
    .reset(PE_11_reset),
    .io_data_2_in_valid(PE_11_io_data_2_in_valid),
    .io_data_2_in_bits(PE_11_io_data_2_in_bits),
    .io_data_2_out_valid(PE_11_io_data_2_out_valid),
    .io_data_2_out_bits(PE_11_io_data_2_out_bits),
    .io_data_1_in_valid(PE_11_io_data_1_in_valid),
    .io_data_1_in_bits(PE_11_io_data_1_in_bits),
    .io_data_1_out_valid(PE_11_io_data_1_out_valid),
    .io_data_1_out_bits(PE_11_io_data_1_out_bits),
    .io_data_0_in_valid(PE_11_io_data_0_in_valid),
    .io_data_0_in_bits(PE_11_io_data_0_in_bits),
    .io_data_0_out_valid(PE_11_io_data_0_out_valid),
    .io_data_0_out_bits(PE_11_io_data_0_out_bits),
    .io_sig_stat2trans(PE_11_io_sig_stat2trans)
  );
  PE PE_12 ( // @[pearray.scala 103:13]
    .clock(PE_12_clock),
    .reset(PE_12_reset),
    .io_data_2_in_valid(PE_12_io_data_2_in_valid),
    .io_data_2_in_bits(PE_12_io_data_2_in_bits),
    .io_data_2_out_valid(PE_12_io_data_2_out_valid),
    .io_data_2_out_bits(PE_12_io_data_2_out_bits),
    .io_data_1_in_valid(PE_12_io_data_1_in_valid),
    .io_data_1_in_bits(PE_12_io_data_1_in_bits),
    .io_data_1_out_valid(PE_12_io_data_1_out_valid),
    .io_data_1_out_bits(PE_12_io_data_1_out_bits),
    .io_data_0_in_valid(PE_12_io_data_0_in_valid),
    .io_data_0_in_bits(PE_12_io_data_0_in_bits),
    .io_data_0_out_valid(PE_12_io_data_0_out_valid),
    .io_data_0_out_bits(PE_12_io_data_0_out_bits),
    .io_sig_stat2trans(PE_12_io_sig_stat2trans)
  );
  PE PE_13 ( // @[pearray.scala 103:13]
    .clock(PE_13_clock),
    .reset(PE_13_reset),
    .io_data_2_in_valid(PE_13_io_data_2_in_valid),
    .io_data_2_in_bits(PE_13_io_data_2_in_bits),
    .io_data_2_out_valid(PE_13_io_data_2_out_valid),
    .io_data_2_out_bits(PE_13_io_data_2_out_bits),
    .io_data_1_in_valid(PE_13_io_data_1_in_valid),
    .io_data_1_in_bits(PE_13_io_data_1_in_bits),
    .io_data_1_out_valid(PE_13_io_data_1_out_valid),
    .io_data_1_out_bits(PE_13_io_data_1_out_bits),
    .io_data_0_in_valid(PE_13_io_data_0_in_valid),
    .io_data_0_in_bits(PE_13_io_data_0_in_bits),
    .io_data_0_out_valid(PE_13_io_data_0_out_valid),
    .io_data_0_out_bits(PE_13_io_data_0_out_bits),
    .io_sig_stat2trans(PE_13_io_sig_stat2trans)
  );
  PE PE_14 ( // @[pearray.scala 103:13]
    .clock(PE_14_clock),
    .reset(PE_14_reset),
    .io_data_2_in_valid(PE_14_io_data_2_in_valid),
    .io_data_2_in_bits(PE_14_io_data_2_in_bits),
    .io_data_2_out_valid(PE_14_io_data_2_out_valid),
    .io_data_2_out_bits(PE_14_io_data_2_out_bits),
    .io_data_1_in_valid(PE_14_io_data_1_in_valid),
    .io_data_1_in_bits(PE_14_io_data_1_in_bits),
    .io_data_1_out_valid(PE_14_io_data_1_out_valid),
    .io_data_1_out_bits(PE_14_io_data_1_out_bits),
    .io_data_0_in_valid(PE_14_io_data_0_in_valid),
    .io_data_0_in_bits(PE_14_io_data_0_in_bits),
    .io_data_0_out_valid(PE_14_io_data_0_out_valid),
    .io_data_0_out_bits(PE_14_io_data_0_out_bits),
    .io_sig_stat2trans(PE_14_io_sig_stat2trans)
  );
  PE PE_15 ( // @[pearray.scala 103:13]
    .clock(PE_15_clock),
    .reset(PE_15_reset),
    .io_data_2_in_valid(PE_15_io_data_2_in_valid),
    .io_data_2_in_bits(PE_15_io_data_2_in_bits),
    .io_data_2_out_valid(PE_15_io_data_2_out_valid),
    .io_data_2_out_bits(PE_15_io_data_2_out_bits),
    .io_data_1_in_valid(PE_15_io_data_1_in_valid),
    .io_data_1_in_bits(PE_15_io_data_1_in_bits),
    .io_data_1_out_valid(PE_15_io_data_1_out_valid),
    .io_data_1_out_bits(PE_15_io_data_1_out_bits),
    .io_data_0_in_valid(PE_15_io_data_0_in_valid),
    .io_data_0_in_bits(PE_15_io_data_0_in_bits),
    .io_data_0_out_valid(PE_15_io_data_0_out_valid),
    .io_data_0_out_bits(PE_15_io_data_0_out_bits),
    .io_sig_stat2trans(PE_15_io_sig_stat2trans)
  );
  PE PE_16 ( // @[pearray.scala 103:13]
    .clock(PE_16_clock),
    .reset(PE_16_reset),
    .io_data_2_in_valid(PE_16_io_data_2_in_valid),
    .io_data_2_in_bits(PE_16_io_data_2_in_bits),
    .io_data_2_out_valid(PE_16_io_data_2_out_valid),
    .io_data_2_out_bits(PE_16_io_data_2_out_bits),
    .io_data_1_in_valid(PE_16_io_data_1_in_valid),
    .io_data_1_in_bits(PE_16_io_data_1_in_bits),
    .io_data_1_out_valid(PE_16_io_data_1_out_valid),
    .io_data_1_out_bits(PE_16_io_data_1_out_bits),
    .io_data_0_in_valid(PE_16_io_data_0_in_valid),
    .io_data_0_in_bits(PE_16_io_data_0_in_bits),
    .io_data_0_out_valid(PE_16_io_data_0_out_valid),
    .io_data_0_out_bits(PE_16_io_data_0_out_bits),
    .io_sig_stat2trans(PE_16_io_sig_stat2trans)
  );
  PE PE_17 ( // @[pearray.scala 103:13]
    .clock(PE_17_clock),
    .reset(PE_17_reset),
    .io_data_2_in_valid(PE_17_io_data_2_in_valid),
    .io_data_2_in_bits(PE_17_io_data_2_in_bits),
    .io_data_2_out_valid(PE_17_io_data_2_out_valid),
    .io_data_2_out_bits(PE_17_io_data_2_out_bits),
    .io_data_1_in_valid(PE_17_io_data_1_in_valid),
    .io_data_1_in_bits(PE_17_io_data_1_in_bits),
    .io_data_1_out_valid(PE_17_io_data_1_out_valid),
    .io_data_1_out_bits(PE_17_io_data_1_out_bits),
    .io_data_0_in_valid(PE_17_io_data_0_in_valid),
    .io_data_0_in_bits(PE_17_io_data_0_in_bits),
    .io_data_0_out_valid(PE_17_io_data_0_out_valid),
    .io_data_0_out_bits(PE_17_io_data_0_out_bits),
    .io_sig_stat2trans(PE_17_io_sig_stat2trans)
  );
  PE PE_18 ( // @[pearray.scala 103:13]
    .clock(PE_18_clock),
    .reset(PE_18_reset),
    .io_data_2_in_valid(PE_18_io_data_2_in_valid),
    .io_data_2_in_bits(PE_18_io_data_2_in_bits),
    .io_data_2_out_valid(PE_18_io_data_2_out_valid),
    .io_data_2_out_bits(PE_18_io_data_2_out_bits),
    .io_data_1_in_valid(PE_18_io_data_1_in_valid),
    .io_data_1_in_bits(PE_18_io_data_1_in_bits),
    .io_data_1_out_valid(PE_18_io_data_1_out_valid),
    .io_data_1_out_bits(PE_18_io_data_1_out_bits),
    .io_data_0_in_valid(PE_18_io_data_0_in_valid),
    .io_data_0_in_bits(PE_18_io_data_0_in_bits),
    .io_data_0_out_valid(PE_18_io_data_0_out_valid),
    .io_data_0_out_bits(PE_18_io_data_0_out_bits),
    .io_sig_stat2trans(PE_18_io_sig_stat2trans)
  );
  PE PE_19 ( // @[pearray.scala 103:13]
    .clock(PE_19_clock),
    .reset(PE_19_reset),
    .io_data_2_in_valid(PE_19_io_data_2_in_valid),
    .io_data_2_in_bits(PE_19_io_data_2_in_bits),
    .io_data_2_out_valid(PE_19_io_data_2_out_valid),
    .io_data_2_out_bits(PE_19_io_data_2_out_bits),
    .io_data_1_in_valid(PE_19_io_data_1_in_valid),
    .io_data_1_in_bits(PE_19_io_data_1_in_bits),
    .io_data_1_out_valid(PE_19_io_data_1_out_valid),
    .io_data_1_out_bits(PE_19_io_data_1_out_bits),
    .io_data_0_in_valid(PE_19_io_data_0_in_valid),
    .io_data_0_in_bits(PE_19_io_data_0_in_bits),
    .io_data_0_out_valid(PE_19_io_data_0_out_valid),
    .io_data_0_out_bits(PE_19_io_data_0_out_bits),
    .io_sig_stat2trans(PE_19_io_sig_stat2trans)
  );
  PE PE_20 ( // @[pearray.scala 103:13]
    .clock(PE_20_clock),
    .reset(PE_20_reset),
    .io_data_2_in_valid(PE_20_io_data_2_in_valid),
    .io_data_2_in_bits(PE_20_io_data_2_in_bits),
    .io_data_2_out_valid(PE_20_io_data_2_out_valid),
    .io_data_2_out_bits(PE_20_io_data_2_out_bits),
    .io_data_1_in_valid(PE_20_io_data_1_in_valid),
    .io_data_1_in_bits(PE_20_io_data_1_in_bits),
    .io_data_1_out_valid(PE_20_io_data_1_out_valid),
    .io_data_1_out_bits(PE_20_io_data_1_out_bits),
    .io_data_0_in_valid(PE_20_io_data_0_in_valid),
    .io_data_0_in_bits(PE_20_io_data_0_in_bits),
    .io_data_0_out_valid(PE_20_io_data_0_out_valid),
    .io_data_0_out_bits(PE_20_io_data_0_out_bits),
    .io_sig_stat2trans(PE_20_io_sig_stat2trans)
  );
  PE PE_21 ( // @[pearray.scala 103:13]
    .clock(PE_21_clock),
    .reset(PE_21_reset),
    .io_data_2_in_valid(PE_21_io_data_2_in_valid),
    .io_data_2_in_bits(PE_21_io_data_2_in_bits),
    .io_data_2_out_valid(PE_21_io_data_2_out_valid),
    .io_data_2_out_bits(PE_21_io_data_2_out_bits),
    .io_data_1_in_valid(PE_21_io_data_1_in_valid),
    .io_data_1_in_bits(PE_21_io_data_1_in_bits),
    .io_data_1_out_valid(PE_21_io_data_1_out_valid),
    .io_data_1_out_bits(PE_21_io_data_1_out_bits),
    .io_data_0_in_valid(PE_21_io_data_0_in_valid),
    .io_data_0_in_bits(PE_21_io_data_0_in_bits),
    .io_data_0_out_valid(PE_21_io_data_0_out_valid),
    .io_data_0_out_bits(PE_21_io_data_0_out_bits),
    .io_sig_stat2trans(PE_21_io_sig_stat2trans)
  );
  PE PE_22 ( // @[pearray.scala 103:13]
    .clock(PE_22_clock),
    .reset(PE_22_reset),
    .io_data_2_in_valid(PE_22_io_data_2_in_valid),
    .io_data_2_in_bits(PE_22_io_data_2_in_bits),
    .io_data_2_out_valid(PE_22_io_data_2_out_valid),
    .io_data_2_out_bits(PE_22_io_data_2_out_bits),
    .io_data_1_in_valid(PE_22_io_data_1_in_valid),
    .io_data_1_in_bits(PE_22_io_data_1_in_bits),
    .io_data_1_out_valid(PE_22_io_data_1_out_valid),
    .io_data_1_out_bits(PE_22_io_data_1_out_bits),
    .io_data_0_in_valid(PE_22_io_data_0_in_valid),
    .io_data_0_in_bits(PE_22_io_data_0_in_bits),
    .io_data_0_out_valid(PE_22_io_data_0_out_valid),
    .io_data_0_out_bits(PE_22_io_data_0_out_bits),
    .io_sig_stat2trans(PE_22_io_sig_stat2trans)
  );
  PE PE_23 ( // @[pearray.scala 103:13]
    .clock(PE_23_clock),
    .reset(PE_23_reset),
    .io_data_2_in_valid(PE_23_io_data_2_in_valid),
    .io_data_2_in_bits(PE_23_io_data_2_in_bits),
    .io_data_2_out_valid(PE_23_io_data_2_out_valid),
    .io_data_2_out_bits(PE_23_io_data_2_out_bits),
    .io_data_1_in_valid(PE_23_io_data_1_in_valid),
    .io_data_1_in_bits(PE_23_io_data_1_in_bits),
    .io_data_1_out_valid(PE_23_io_data_1_out_valid),
    .io_data_1_out_bits(PE_23_io_data_1_out_bits),
    .io_data_0_in_valid(PE_23_io_data_0_in_valid),
    .io_data_0_in_bits(PE_23_io_data_0_in_bits),
    .io_data_0_out_valid(PE_23_io_data_0_out_valid),
    .io_data_0_out_bits(PE_23_io_data_0_out_bits),
    .io_sig_stat2trans(PE_23_io_sig_stat2trans)
  );
  PE PE_24 ( // @[pearray.scala 103:13]
    .clock(PE_24_clock),
    .reset(PE_24_reset),
    .io_data_2_in_valid(PE_24_io_data_2_in_valid),
    .io_data_2_in_bits(PE_24_io_data_2_in_bits),
    .io_data_2_out_valid(PE_24_io_data_2_out_valid),
    .io_data_2_out_bits(PE_24_io_data_2_out_bits),
    .io_data_1_in_valid(PE_24_io_data_1_in_valid),
    .io_data_1_in_bits(PE_24_io_data_1_in_bits),
    .io_data_1_out_valid(PE_24_io_data_1_out_valid),
    .io_data_1_out_bits(PE_24_io_data_1_out_bits),
    .io_data_0_in_valid(PE_24_io_data_0_in_valid),
    .io_data_0_in_bits(PE_24_io_data_0_in_bits),
    .io_data_0_out_valid(PE_24_io_data_0_out_valid),
    .io_data_0_out_bits(PE_24_io_data_0_out_bits),
    .io_sig_stat2trans(PE_24_io_sig_stat2trans)
  );
  PE PE_25 ( // @[pearray.scala 103:13]
    .clock(PE_25_clock),
    .reset(PE_25_reset),
    .io_data_2_in_valid(PE_25_io_data_2_in_valid),
    .io_data_2_in_bits(PE_25_io_data_2_in_bits),
    .io_data_2_out_valid(PE_25_io_data_2_out_valid),
    .io_data_2_out_bits(PE_25_io_data_2_out_bits),
    .io_data_1_in_valid(PE_25_io_data_1_in_valid),
    .io_data_1_in_bits(PE_25_io_data_1_in_bits),
    .io_data_1_out_valid(PE_25_io_data_1_out_valid),
    .io_data_1_out_bits(PE_25_io_data_1_out_bits),
    .io_data_0_in_valid(PE_25_io_data_0_in_valid),
    .io_data_0_in_bits(PE_25_io_data_0_in_bits),
    .io_data_0_out_valid(PE_25_io_data_0_out_valid),
    .io_data_0_out_bits(PE_25_io_data_0_out_bits),
    .io_sig_stat2trans(PE_25_io_sig_stat2trans)
  );
  PE PE_26 ( // @[pearray.scala 103:13]
    .clock(PE_26_clock),
    .reset(PE_26_reset),
    .io_data_2_in_valid(PE_26_io_data_2_in_valid),
    .io_data_2_in_bits(PE_26_io_data_2_in_bits),
    .io_data_2_out_valid(PE_26_io_data_2_out_valid),
    .io_data_2_out_bits(PE_26_io_data_2_out_bits),
    .io_data_1_in_valid(PE_26_io_data_1_in_valid),
    .io_data_1_in_bits(PE_26_io_data_1_in_bits),
    .io_data_1_out_valid(PE_26_io_data_1_out_valid),
    .io_data_1_out_bits(PE_26_io_data_1_out_bits),
    .io_data_0_in_valid(PE_26_io_data_0_in_valid),
    .io_data_0_in_bits(PE_26_io_data_0_in_bits),
    .io_data_0_out_valid(PE_26_io_data_0_out_valid),
    .io_data_0_out_bits(PE_26_io_data_0_out_bits),
    .io_sig_stat2trans(PE_26_io_sig_stat2trans)
  );
  PE PE_27 ( // @[pearray.scala 103:13]
    .clock(PE_27_clock),
    .reset(PE_27_reset),
    .io_data_2_in_valid(PE_27_io_data_2_in_valid),
    .io_data_2_in_bits(PE_27_io_data_2_in_bits),
    .io_data_2_out_valid(PE_27_io_data_2_out_valid),
    .io_data_2_out_bits(PE_27_io_data_2_out_bits),
    .io_data_1_in_valid(PE_27_io_data_1_in_valid),
    .io_data_1_in_bits(PE_27_io_data_1_in_bits),
    .io_data_1_out_valid(PE_27_io_data_1_out_valid),
    .io_data_1_out_bits(PE_27_io_data_1_out_bits),
    .io_data_0_in_valid(PE_27_io_data_0_in_valid),
    .io_data_0_in_bits(PE_27_io_data_0_in_bits),
    .io_data_0_out_valid(PE_27_io_data_0_out_valid),
    .io_data_0_out_bits(PE_27_io_data_0_out_bits),
    .io_sig_stat2trans(PE_27_io_sig_stat2trans)
  );
  PE PE_28 ( // @[pearray.scala 103:13]
    .clock(PE_28_clock),
    .reset(PE_28_reset),
    .io_data_2_in_valid(PE_28_io_data_2_in_valid),
    .io_data_2_in_bits(PE_28_io_data_2_in_bits),
    .io_data_2_out_valid(PE_28_io_data_2_out_valid),
    .io_data_2_out_bits(PE_28_io_data_2_out_bits),
    .io_data_1_in_valid(PE_28_io_data_1_in_valid),
    .io_data_1_in_bits(PE_28_io_data_1_in_bits),
    .io_data_1_out_valid(PE_28_io_data_1_out_valid),
    .io_data_1_out_bits(PE_28_io_data_1_out_bits),
    .io_data_0_in_valid(PE_28_io_data_0_in_valid),
    .io_data_0_in_bits(PE_28_io_data_0_in_bits),
    .io_data_0_out_valid(PE_28_io_data_0_out_valid),
    .io_data_0_out_bits(PE_28_io_data_0_out_bits),
    .io_sig_stat2trans(PE_28_io_sig_stat2trans)
  );
  PE PE_29 ( // @[pearray.scala 103:13]
    .clock(PE_29_clock),
    .reset(PE_29_reset),
    .io_data_2_in_valid(PE_29_io_data_2_in_valid),
    .io_data_2_in_bits(PE_29_io_data_2_in_bits),
    .io_data_2_out_valid(PE_29_io_data_2_out_valid),
    .io_data_2_out_bits(PE_29_io_data_2_out_bits),
    .io_data_1_in_valid(PE_29_io_data_1_in_valid),
    .io_data_1_in_bits(PE_29_io_data_1_in_bits),
    .io_data_1_out_valid(PE_29_io_data_1_out_valid),
    .io_data_1_out_bits(PE_29_io_data_1_out_bits),
    .io_data_0_in_valid(PE_29_io_data_0_in_valid),
    .io_data_0_in_bits(PE_29_io_data_0_in_bits),
    .io_data_0_out_valid(PE_29_io_data_0_out_valid),
    .io_data_0_out_bits(PE_29_io_data_0_out_bits),
    .io_sig_stat2trans(PE_29_io_sig_stat2trans)
  );
  PE PE_30 ( // @[pearray.scala 103:13]
    .clock(PE_30_clock),
    .reset(PE_30_reset),
    .io_data_2_in_valid(PE_30_io_data_2_in_valid),
    .io_data_2_in_bits(PE_30_io_data_2_in_bits),
    .io_data_2_out_valid(PE_30_io_data_2_out_valid),
    .io_data_2_out_bits(PE_30_io_data_2_out_bits),
    .io_data_1_in_valid(PE_30_io_data_1_in_valid),
    .io_data_1_in_bits(PE_30_io_data_1_in_bits),
    .io_data_1_out_valid(PE_30_io_data_1_out_valid),
    .io_data_1_out_bits(PE_30_io_data_1_out_bits),
    .io_data_0_in_valid(PE_30_io_data_0_in_valid),
    .io_data_0_in_bits(PE_30_io_data_0_in_bits),
    .io_data_0_out_valid(PE_30_io_data_0_out_valid),
    .io_data_0_out_bits(PE_30_io_data_0_out_bits),
    .io_sig_stat2trans(PE_30_io_sig_stat2trans)
  );
  PE PE_31 ( // @[pearray.scala 103:13]
    .clock(PE_31_clock),
    .reset(PE_31_reset),
    .io_data_2_in_valid(PE_31_io_data_2_in_valid),
    .io_data_2_in_bits(PE_31_io_data_2_in_bits),
    .io_data_2_out_valid(PE_31_io_data_2_out_valid),
    .io_data_2_out_bits(PE_31_io_data_2_out_bits),
    .io_data_1_in_valid(PE_31_io_data_1_in_valid),
    .io_data_1_in_bits(PE_31_io_data_1_in_bits),
    .io_data_1_out_valid(PE_31_io_data_1_out_valid),
    .io_data_1_out_bits(PE_31_io_data_1_out_bits),
    .io_data_0_in_valid(PE_31_io_data_0_in_valid),
    .io_data_0_in_bits(PE_31_io_data_0_in_bits),
    .io_data_0_out_valid(PE_31_io_data_0_out_valid),
    .io_data_0_out_bits(PE_31_io_data_0_out_bits),
    .io_sig_stat2trans(PE_31_io_sig_stat2trans)
  );
  PE PE_32 ( // @[pearray.scala 103:13]
    .clock(PE_32_clock),
    .reset(PE_32_reset),
    .io_data_2_in_valid(PE_32_io_data_2_in_valid),
    .io_data_2_in_bits(PE_32_io_data_2_in_bits),
    .io_data_2_out_valid(PE_32_io_data_2_out_valid),
    .io_data_2_out_bits(PE_32_io_data_2_out_bits),
    .io_data_1_in_valid(PE_32_io_data_1_in_valid),
    .io_data_1_in_bits(PE_32_io_data_1_in_bits),
    .io_data_1_out_valid(PE_32_io_data_1_out_valid),
    .io_data_1_out_bits(PE_32_io_data_1_out_bits),
    .io_data_0_in_valid(PE_32_io_data_0_in_valid),
    .io_data_0_in_bits(PE_32_io_data_0_in_bits),
    .io_data_0_out_valid(PE_32_io_data_0_out_valid),
    .io_data_0_out_bits(PE_32_io_data_0_out_bits),
    .io_sig_stat2trans(PE_32_io_sig_stat2trans)
  );
  PE PE_33 ( // @[pearray.scala 103:13]
    .clock(PE_33_clock),
    .reset(PE_33_reset),
    .io_data_2_in_valid(PE_33_io_data_2_in_valid),
    .io_data_2_in_bits(PE_33_io_data_2_in_bits),
    .io_data_2_out_valid(PE_33_io_data_2_out_valid),
    .io_data_2_out_bits(PE_33_io_data_2_out_bits),
    .io_data_1_in_valid(PE_33_io_data_1_in_valid),
    .io_data_1_in_bits(PE_33_io_data_1_in_bits),
    .io_data_1_out_valid(PE_33_io_data_1_out_valid),
    .io_data_1_out_bits(PE_33_io_data_1_out_bits),
    .io_data_0_in_valid(PE_33_io_data_0_in_valid),
    .io_data_0_in_bits(PE_33_io_data_0_in_bits),
    .io_data_0_out_valid(PE_33_io_data_0_out_valid),
    .io_data_0_out_bits(PE_33_io_data_0_out_bits),
    .io_sig_stat2trans(PE_33_io_sig_stat2trans)
  );
  PE PE_34 ( // @[pearray.scala 103:13]
    .clock(PE_34_clock),
    .reset(PE_34_reset),
    .io_data_2_in_valid(PE_34_io_data_2_in_valid),
    .io_data_2_in_bits(PE_34_io_data_2_in_bits),
    .io_data_2_out_valid(PE_34_io_data_2_out_valid),
    .io_data_2_out_bits(PE_34_io_data_2_out_bits),
    .io_data_1_in_valid(PE_34_io_data_1_in_valid),
    .io_data_1_in_bits(PE_34_io_data_1_in_bits),
    .io_data_1_out_valid(PE_34_io_data_1_out_valid),
    .io_data_1_out_bits(PE_34_io_data_1_out_bits),
    .io_data_0_in_valid(PE_34_io_data_0_in_valid),
    .io_data_0_in_bits(PE_34_io_data_0_in_bits),
    .io_data_0_out_valid(PE_34_io_data_0_out_valid),
    .io_data_0_out_bits(PE_34_io_data_0_out_bits),
    .io_sig_stat2trans(PE_34_io_sig_stat2trans)
  );
  PE PE_35 ( // @[pearray.scala 103:13]
    .clock(PE_35_clock),
    .reset(PE_35_reset),
    .io_data_2_in_valid(PE_35_io_data_2_in_valid),
    .io_data_2_in_bits(PE_35_io_data_2_in_bits),
    .io_data_2_out_valid(PE_35_io_data_2_out_valid),
    .io_data_2_out_bits(PE_35_io_data_2_out_bits),
    .io_data_1_in_valid(PE_35_io_data_1_in_valid),
    .io_data_1_in_bits(PE_35_io_data_1_in_bits),
    .io_data_1_out_valid(PE_35_io_data_1_out_valid),
    .io_data_1_out_bits(PE_35_io_data_1_out_bits),
    .io_data_0_in_valid(PE_35_io_data_0_in_valid),
    .io_data_0_in_bits(PE_35_io_data_0_in_bits),
    .io_data_0_out_valid(PE_35_io_data_0_out_valid),
    .io_data_0_out_bits(PE_35_io_data_0_out_bits),
    .io_sig_stat2trans(PE_35_io_sig_stat2trans)
  );
  PE PE_36 ( // @[pearray.scala 103:13]
    .clock(PE_36_clock),
    .reset(PE_36_reset),
    .io_data_2_in_valid(PE_36_io_data_2_in_valid),
    .io_data_2_in_bits(PE_36_io_data_2_in_bits),
    .io_data_2_out_valid(PE_36_io_data_2_out_valid),
    .io_data_2_out_bits(PE_36_io_data_2_out_bits),
    .io_data_1_in_valid(PE_36_io_data_1_in_valid),
    .io_data_1_in_bits(PE_36_io_data_1_in_bits),
    .io_data_1_out_valid(PE_36_io_data_1_out_valid),
    .io_data_1_out_bits(PE_36_io_data_1_out_bits),
    .io_data_0_in_valid(PE_36_io_data_0_in_valid),
    .io_data_0_in_bits(PE_36_io_data_0_in_bits),
    .io_data_0_out_valid(PE_36_io_data_0_out_valid),
    .io_data_0_out_bits(PE_36_io_data_0_out_bits),
    .io_sig_stat2trans(PE_36_io_sig_stat2trans)
  );
  PE PE_37 ( // @[pearray.scala 103:13]
    .clock(PE_37_clock),
    .reset(PE_37_reset),
    .io_data_2_in_valid(PE_37_io_data_2_in_valid),
    .io_data_2_in_bits(PE_37_io_data_2_in_bits),
    .io_data_2_out_valid(PE_37_io_data_2_out_valid),
    .io_data_2_out_bits(PE_37_io_data_2_out_bits),
    .io_data_1_in_valid(PE_37_io_data_1_in_valid),
    .io_data_1_in_bits(PE_37_io_data_1_in_bits),
    .io_data_1_out_valid(PE_37_io_data_1_out_valid),
    .io_data_1_out_bits(PE_37_io_data_1_out_bits),
    .io_data_0_in_valid(PE_37_io_data_0_in_valid),
    .io_data_0_in_bits(PE_37_io_data_0_in_bits),
    .io_data_0_out_valid(PE_37_io_data_0_out_valid),
    .io_data_0_out_bits(PE_37_io_data_0_out_bits),
    .io_sig_stat2trans(PE_37_io_sig_stat2trans)
  );
  PE PE_38 ( // @[pearray.scala 103:13]
    .clock(PE_38_clock),
    .reset(PE_38_reset),
    .io_data_2_in_valid(PE_38_io_data_2_in_valid),
    .io_data_2_in_bits(PE_38_io_data_2_in_bits),
    .io_data_2_out_valid(PE_38_io_data_2_out_valid),
    .io_data_2_out_bits(PE_38_io_data_2_out_bits),
    .io_data_1_in_valid(PE_38_io_data_1_in_valid),
    .io_data_1_in_bits(PE_38_io_data_1_in_bits),
    .io_data_1_out_valid(PE_38_io_data_1_out_valid),
    .io_data_1_out_bits(PE_38_io_data_1_out_bits),
    .io_data_0_in_valid(PE_38_io_data_0_in_valid),
    .io_data_0_in_bits(PE_38_io_data_0_in_bits),
    .io_data_0_out_valid(PE_38_io_data_0_out_valid),
    .io_data_0_out_bits(PE_38_io_data_0_out_bits),
    .io_sig_stat2trans(PE_38_io_sig_stat2trans)
  );
  PE PE_39 ( // @[pearray.scala 103:13]
    .clock(PE_39_clock),
    .reset(PE_39_reset),
    .io_data_2_in_valid(PE_39_io_data_2_in_valid),
    .io_data_2_in_bits(PE_39_io_data_2_in_bits),
    .io_data_2_out_valid(PE_39_io_data_2_out_valid),
    .io_data_2_out_bits(PE_39_io_data_2_out_bits),
    .io_data_1_in_valid(PE_39_io_data_1_in_valid),
    .io_data_1_in_bits(PE_39_io_data_1_in_bits),
    .io_data_1_out_valid(PE_39_io_data_1_out_valid),
    .io_data_1_out_bits(PE_39_io_data_1_out_bits),
    .io_data_0_in_valid(PE_39_io_data_0_in_valid),
    .io_data_0_in_bits(PE_39_io_data_0_in_bits),
    .io_data_0_out_valid(PE_39_io_data_0_out_valid),
    .io_data_0_out_bits(PE_39_io_data_0_out_bits),
    .io_sig_stat2trans(PE_39_io_sig_stat2trans)
  );
  PE PE_40 ( // @[pearray.scala 103:13]
    .clock(PE_40_clock),
    .reset(PE_40_reset),
    .io_data_2_in_valid(PE_40_io_data_2_in_valid),
    .io_data_2_in_bits(PE_40_io_data_2_in_bits),
    .io_data_2_out_valid(PE_40_io_data_2_out_valid),
    .io_data_2_out_bits(PE_40_io_data_2_out_bits),
    .io_data_1_in_valid(PE_40_io_data_1_in_valid),
    .io_data_1_in_bits(PE_40_io_data_1_in_bits),
    .io_data_1_out_valid(PE_40_io_data_1_out_valid),
    .io_data_1_out_bits(PE_40_io_data_1_out_bits),
    .io_data_0_in_valid(PE_40_io_data_0_in_valid),
    .io_data_0_in_bits(PE_40_io_data_0_in_bits),
    .io_data_0_out_valid(PE_40_io_data_0_out_valid),
    .io_data_0_out_bits(PE_40_io_data_0_out_bits),
    .io_sig_stat2trans(PE_40_io_sig_stat2trans)
  );
  PE PE_41 ( // @[pearray.scala 103:13]
    .clock(PE_41_clock),
    .reset(PE_41_reset),
    .io_data_2_in_valid(PE_41_io_data_2_in_valid),
    .io_data_2_in_bits(PE_41_io_data_2_in_bits),
    .io_data_2_out_valid(PE_41_io_data_2_out_valid),
    .io_data_2_out_bits(PE_41_io_data_2_out_bits),
    .io_data_1_in_valid(PE_41_io_data_1_in_valid),
    .io_data_1_in_bits(PE_41_io_data_1_in_bits),
    .io_data_1_out_valid(PE_41_io_data_1_out_valid),
    .io_data_1_out_bits(PE_41_io_data_1_out_bits),
    .io_data_0_in_valid(PE_41_io_data_0_in_valid),
    .io_data_0_in_bits(PE_41_io_data_0_in_bits),
    .io_data_0_out_valid(PE_41_io_data_0_out_valid),
    .io_data_0_out_bits(PE_41_io_data_0_out_bits),
    .io_sig_stat2trans(PE_41_io_sig_stat2trans)
  );
  PE PE_42 ( // @[pearray.scala 103:13]
    .clock(PE_42_clock),
    .reset(PE_42_reset),
    .io_data_2_in_valid(PE_42_io_data_2_in_valid),
    .io_data_2_in_bits(PE_42_io_data_2_in_bits),
    .io_data_2_out_valid(PE_42_io_data_2_out_valid),
    .io_data_2_out_bits(PE_42_io_data_2_out_bits),
    .io_data_1_in_valid(PE_42_io_data_1_in_valid),
    .io_data_1_in_bits(PE_42_io_data_1_in_bits),
    .io_data_1_out_valid(PE_42_io_data_1_out_valid),
    .io_data_1_out_bits(PE_42_io_data_1_out_bits),
    .io_data_0_in_valid(PE_42_io_data_0_in_valid),
    .io_data_0_in_bits(PE_42_io_data_0_in_bits),
    .io_data_0_out_valid(PE_42_io_data_0_out_valid),
    .io_data_0_out_bits(PE_42_io_data_0_out_bits),
    .io_sig_stat2trans(PE_42_io_sig_stat2trans)
  );
  PE PE_43 ( // @[pearray.scala 103:13]
    .clock(PE_43_clock),
    .reset(PE_43_reset),
    .io_data_2_in_valid(PE_43_io_data_2_in_valid),
    .io_data_2_in_bits(PE_43_io_data_2_in_bits),
    .io_data_2_out_valid(PE_43_io_data_2_out_valid),
    .io_data_2_out_bits(PE_43_io_data_2_out_bits),
    .io_data_1_in_valid(PE_43_io_data_1_in_valid),
    .io_data_1_in_bits(PE_43_io_data_1_in_bits),
    .io_data_1_out_valid(PE_43_io_data_1_out_valid),
    .io_data_1_out_bits(PE_43_io_data_1_out_bits),
    .io_data_0_in_valid(PE_43_io_data_0_in_valid),
    .io_data_0_in_bits(PE_43_io_data_0_in_bits),
    .io_data_0_out_valid(PE_43_io_data_0_out_valid),
    .io_data_0_out_bits(PE_43_io_data_0_out_bits),
    .io_sig_stat2trans(PE_43_io_sig_stat2trans)
  );
  PE PE_44 ( // @[pearray.scala 103:13]
    .clock(PE_44_clock),
    .reset(PE_44_reset),
    .io_data_2_in_valid(PE_44_io_data_2_in_valid),
    .io_data_2_in_bits(PE_44_io_data_2_in_bits),
    .io_data_2_out_valid(PE_44_io_data_2_out_valid),
    .io_data_2_out_bits(PE_44_io_data_2_out_bits),
    .io_data_1_in_valid(PE_44_io_data_1_in_valid),
    .io_data_1_in_bits(PE_44_io_data_1_in_bits),
    .io_data_1_out_valid(PE_44_io_data_1_out_valid),
    .io_data_1_out_bits(PE_44_io_data_1_out_bits),
    .io_data_0_in_valid(PE_44_io_data_0_in_valid),
    .io_data_0_in_bits(PE_44_io_data_0_in_bits),
    .io_data_0_out_valid(PE_44_io_data_0_out_valid),
    .io_data_0_out_bits(PE_44_io_data_0_out_bits),
    .io_sig_stat2trans(PE_44_io_sig_stat2trans)
  );
  PE PE_45 ( // @[pearray.scala 103:13]
    .clock(PE_45_clock),
    .reset(PE_45_reset),
    .io_data_2_in_valid(PE_45_io_data_2_in_valid),
    .io_data_2_in_bits(PE_45_io_data_2_in_bits),
    .io_data_2_out_valid(PE_45_io_data_2_out_valid),
    .io_data_2_out_bits(PE_45_io_data_2_out_bits),
    .io_data_1_in_valid(PE_45_io_data_1_in_valid),
    .io_data_1_in_bits(PE_45_io_data_1_in_bits),
    .io_data_1_out_valid(PE_45_io_data_1_out_valid),
    .io_data_1_out_bits(PE_45_io_data_1_out_bits),
    .io_data_0_in_valid(PE_45_io_data_0_in_valid),
    .io_data_0_in_bits(PE_45_io_data_0_in_bits),
    .io_data_0_out_valid(PE_45_io_data_0_out_valid),
    .io_data_0_out_bits(PE_45_io_data_0_out_bits),
    .io_sig_stat2trans(PE_45_io_sig_stat2trans)
  );
  PE PE_46 ( // @[pearray.scala 103:13]
    .clock(PE_46_clock),
    .reset(PE_46_reset),
    .io_data_2_in_valid(PE_46_io_data_2_in_valid),
    .io_data_2_in_bits(PE_46_io_data_2_in_bits),
    .io_data_2_out_valid(PE_46_io_data_2_out_valid),
    .io_data_2_out_bits(PE_46_io_data_2_out_bits),
    .io_data_1_in_valid(PE_46_io_data_1_in_valid),
    .io_data_1_in_bits(PE_46_io_data_1_in_bits),
    .io_data_1_out_valid(PE_46_io_data_1_out_valid),
    .io_data_1_out_bits(PE_46_io_data_1_out_bits),
    .io_data_0_in_valid(PE_46_io_data_0_in_valid),
    .io_data_0_in_bits(PE_46_io_data_0_in_bits),
    .io_data_0_out_valid(PE_46_io_data_0_out_valid),
    .io_data_0_out_bits(PE_46_io_data_0_out_bits),
    .io_sig_stat2trans(PE_46_io_sig_stat2trans)
  );
  PE PE_47 ( // @[pearray.scala 103:13]
    .clock(PE_47_clock),
    .reset(PE_47_reset),
    .io_data_2_in_valid(PE_47_io_data_2_in_valid),
    .io_data_2_in_bits(PE_47_io_data_2_in_bits),
    .io_data_2_out_valid(PE_47_io_data_2_out_valid),
    .io_data_2_out_bits(PE_47_io_data_2_out_bits),
    .io_data_1_in_valid(PE_47_io_data_1_in_valid),
    .io_data_1_in_bits(PE_47_io_data_1_in_bits),
    .io_data_1_out_valid(PE_47_io_data_1_out_valid),
    .io_data_1_out_bits(PE_47_io_data_1_out_bits),
    .io_data_0_in_valid(PE_47_io_data_0_in_valid),
    .io_data_0_in_bits(PE_47_io_data_0_in_bits),
    .io_data_0_out_valid(PE_47_io_data_0_out_valid),
    .io_data_0_out_bits(PE_47_io_data_0_out_bits),
    .io_sig_stat2trans(PE_47_io_sig_stat2trans)
  );
  PE PE_48 ( // @[pearray.scala 103:13]
    .clock(PE_48_clock),
    .reset(PE_48_reset),
    .io_data_2_in_valid(PE_48_io_data_2_in_valid),
    .io_data_2_in_bits(PE_48_io_data_2_in_bits),
    .io_data_2_out_valid(PE_48_io_data_2_out_valid),
    .io_data_2_out_bits(PE_48_io_data_2_out_bits),
    .io_data_1_in_valid(PE_48_io_data_1_in_valid),
    .io_data_1_in_bits(PE_48_io_data_1_in_bits),
    .io_data_1_out_valid(PE_48_io_data_1_out_valid),
    .io_data_1_out_bits(PE_48_io_data_1_out_bits),
    .io_data_0_in_valid(PE_48_io_data_0_in_valid),
    .io_data_0_in_bits(PE_48_io_data_0_in_bits),
    .io_data_0_out_valid(PE_48_io_data_0_out_valid),
    .io_data_0_out_bits(PE_48_io_data_0_out_bits),
    .io_sig_stat2trans(PE_48_io_sig_stat2trans)
  );
  PE PE_49 ( // @[pearray.scala 103:13]
    .clock(PE_49_clock),
    .reset(PE_49_reset),
    .io_data_2_in_valid(PE_49_io_data_2_in_valid),
    .io_data_2_in_bits(PE_49_io_data_2_in_bits),
    .io_data_2_out_valid(PE_49_io_data_2_out_valid),
    .io_data_2_out_bits(PE_49_io_data_2_out_bits),
    .io_data_1_in_valid(PE_49_io_data_1_in_valid),
    .io_data_1_in_bits(PE_49_io_data_1_in_bits),
    .io_data_1_out_valid(PE_49_io_data_1_out_valid),
    .io_data_1_out_bits(PE_49_io_data_1_out_bits),
    .io_data_0_in_valid(PE_49_io_data_0_in_valid),
    .io_data_0_in_bits(PE_49_io_data_0_in_bits),
    .io_data_0_out_valid(PE_49_io_data_0_out_valid),
    .io_data_0_out_bits(PE_49_io_data_0_out_bits),
    .io_sig_stat2trans(PE_49_io_sig_stat2trans)
  );
  PE PE_50 ( // @[pearray.scala 103:13]
    .clock(PE_50_clock),
    .reset(PE_50_reset),
    .io_data_2_in_valid(PE_50_io_data_2_in_valid),
    .io_data_2_in_bits(PE_50_io_data_2_in_bits),
    .io_data_2_out_valid(PE_50_io_data_2_out_valid),
    .io_data_2_out_bits(PE_50_io_data_2_out_bits),
    .io_data_1_in_valid(PE_50_io_data_1_in_valid),
    .io_data_1_in_bits(PE_50_io_data_1_in_bits),
    .io_data_1_out_valid(PE_50_io_data_1_out_valid),
    .io_data_1_out_bits(PE_50_io_data_1_out_bits),
    .io_data_0_in_valid(PE_50_io_data_0_in_valid),
    .io_data_0_in_bits(PE_50_io_data_0_in_bits),
    .io_data_0_out_valid(PE_50_io_data_0_out_valid),
    .io_data_0_out_bits(PE_50_io_data_0_out_bits),
    .io_sig_stat2trans(PE_50_io_sig_stat2trans)
  );
  PE PE_51 ( // @[pearray.scala 103:13]
    .clock(PE_51_clock),
    .reset(PE_51_reset),
    .io_data_2_in_valid(PE_51_io_data_2_in_valid),
    .io_data_2_in_bits(PE_51_io_data_2_in_bits),
    .io_data_2_out_valid(PE_51_io_data_2_out_valid),
    .io_data_2_out_bits(PE_51_io_data_2_out_bits),
    .io_data_1_in_valid(PE_51_io_data_1_in_valid),
    .io_data_1_in_bits(PE_51_io_data_1_in_bits),
    .io_data_1_out_valid(PE_51_io_data_1_out_valid),
    .io_data_1_out_bits(PE_51_io_data_1_out_bits),
    .io_data_0_in_valid(PE_51_io_data_0_in_valid),
    .io_data_0_in_bits(PE_51_io_data_0_in_bits),
    .io_data_0_out_valid(PE_51_io_data_0_out_valid),
    .io_data_0_out_bits(PE_51_io_data_0_out_bits),
    .io_sig_stat2trans(PE_51_io_sig_stat2trans)
  );
  PE PE_52 ( // @[pearray.scala 103:13]
    .clock(PE_52_clock),
    .reset(PE_52_reset),
    .io_data_2_in_valid(PE_52_io_data_2_in_valid),
    .io_data_2_in_bits(PE_52_io_data_2_in_bits),
    .io_data_2_out_valid(PE_52_io_data_2_out_valid),
    .io_data_2_out_bits(PE_52_io_data_2_out_bits),
    .io_data_1_in_valid(PE_52_io_data_1_in_valid),
    .io_data_1_in_bits(PE_52_io_data_1_in_bits),
    .io_data_1_out_valid(PE_52_io_data_1_out_valid),
    .io_data_1_out_bits(PE_52_io_data_1_out_bits),
    .io_data_0_in_valid(PE_52_io_data_0_in_valid),
    .io_data_0_in_bits(PE_52_io_data_0_in_bits),
    .io_data_0_out_valid(PE_52_io_data_0_out_valid),
    .io_data_0_out_bits(PE_52_io_data_0_out_bits),
    .io_sig_stat2trans(PE_52_io_sig_stat2trans)
  );
  PE PE_53 ( // @[pearray.scala 103:13]
    .clock(PE_53_clock),
    .reset(PE_53_reset),
    .io_data_2_in_valid(PE_53_io_data_2_in_valid),
    .io_data_2_in_bits(PE_53_io_data_2_in_bits),
    .io_data_2_out_valid(PE_53_io_data_2_out_valid),
    .io_data_2_out_bits(PE_53_io_data_2_out_bits),
    .io_data_1_in_valid(PE_53_io_data_1_in_valid),
    .io_data_1_in_bits(PE_53_io_data_1_in_bits),
    .io_data_1_out_valid(PE_53_io_data_1_out_valid),
    .io_data_1_out_bits(PE_53_io_data_1_out_bits),
    .io_data_0_in_valid(PE_53_io_data_0_in_valid),
    .io_data_0_in_bits(PE_53_io_data_0_in_bits),
    .io_data_0_out_valid(PE_53_io_data_0_out_valid),
    .io_data_0_out_bits(PE_53_io_data_0_out_bits),
    .io_sig_stat2trans(PE_53_io_sig_stat2trans)
  );
  PE PE_54 ( // @[pearray.scala 103:13]
    .clock(PE_54_clock),
    .reset(PE_54_reset),
    .io_data_2_in_valid(PE_54_io_data_2_in_valid),
    .io_data_2_in_bits(PE_54_io_data_2_in_bits),
    .io_data_2_out_valid(PE_54_io_data_2_out_valid),
    .io_data_2_out_bits(PE_54_io_data_2_out_bits),
    .io_data_1_in_valid(PE_54_io_data_1_in_valid),
    .io_data_1_in_bits(PE_54_io_data_1_in_bits),
    .io_data_1_out_valid(PE_54_io_data_1_out_valid),
    .io_data_1_out_bits(PE_54_io_data_1_out_bits),
    .io_data_0_in_valid(PE_54_io_data_0_in_valid),
    .io_data_0_in_bits(PE_54_io_data_0_in_bits),
    .io_data_0_out_valid(PE_54_io_data_0_out_valid),
    .io_data_0_out_bits(PE_54_io_data_0_out_bits),
    .io_sig_stat2trans(PE_54_io_sig_stat2trans)
  );
  PE PE_55 ( // @[pearray.scala 103:13]
    .clock(PE_55_clock),
    .reset(PE_55_reset),
    .io_data_2_in_valid(PE_55_io_data_2_in_valid),
    .io_data_2_in_bits(PE_55_io_data_2_in_bits),
    .io_data_2_out_valid(PE_55_io_data_2_out_valid),
    .io_data_2_out_bits(PE_55_io_data_2_out_bits),
    .io_data_1_in_valid(PE_55_io_data_1_in_valid),
    .io_data_1_in_bits(PE_55_io_data_1_in_bits),
    .io_data_1_out_valid(PE_55_io_data_1_out_valid),
    .io_data_1_out_bits(PE_55_io_data_1_out_bits),
    .io_data_0_in_valid(PE_55_io_data_0_in_valid),
    .io_data_0_in_bits(PE_55_io_data_0_in_bits),
    .io_data_0_out_valid(PE_55_io_data_0_out_valid),
    .io_data_0_out_bits(PE_55_io_data_0_out_bits),
    .io_sig_stat2trans(PE_55_io_sig_stat2trans)
  );
  PE PE_56 ( // @[pearray.scala 103:13]
    .clock(PE_56_clock),
    .reset(PE_56_reset),
    .io_data_2_in_valid(PE_56_io_data_2_in_valid),
    .io_data_2_in_bits(PE_56_io_data_2_in_bits),
    .io_data_2_out_valid(PE_56_io_data_2_out_valid),
    .io_data_2_out_bits(PE_56_io_data_2_out_bits),
    .io_data_1_in_valid(PE_56_io_data_1_in_valid),
    .io_data_1_in_bits(PE_56_io_data_1_in_bits),
    .io_data_1_out_valid(PE_56_io_data_1_out_valid),
    .io_data_1_out_bits(PE_56_io_data_1_out_bits),
    .io_data_0_in_valid(PE_56_io_data_0_in_valid),
    .io_data_0_in_bits(PE_56_io_data_0_in_bits),
    .io_data_0_out_valid(PE_56_io_data_0_out_valid),
    .io_data_0_out_bits(PE_56_io_data_0_out_bits),
    .io_sig_stat2trans(PE_56_io_sig_stat2trans)
  );
  PE PE_57 ( // @[pearray.scala 103:13]
    .clock(PE_57_clock),
    .reset(PE_57_reset),
    .io_data_2_in_valid(PE_57_io_data_2_in_valid),
    .io_data_2_in_bits(PE_57_io_data_2_in_bits),
    .io_data_2_out_valid(PE_57_io_data_2_out_valid),
    .io_data_2_out_bits(PE_57_io_data_2_out_bits),
    .io_data_1_in_valid(PE_57_io_data_1_in_valid),
    .io_data_1_in_bits(PE_57_io_data_1_in_bits),
    .io_data_1_out_valid(PE_57_io_data_1_out_valid),
    .io_data_1_out_bits(PE_57_io_data_1_out_bits),
    .io_data_0_in_valid(PE_57_io_data_0_in_valid),
    .io_data_0_in_bits(PE_57_io_data_0_in_bits),
    .io_data_0_out_valid(PE_57_io_data_0_out_valid),
    .io_data_0_out_bits(PE_57_io_data_0_out_bits),
    .io_sig_stat2trans(PE_57_io_sig_stat2trans)
  );
  PE PE_58 ( // @[pearray.scala 103:13]
    .clock(PE_58_clock),
    .reset(PE_58_reset),
    .io_data_2_in_valid(PE_58_io_data_2_in_valid),
    .io_data_2_in_bits(PE_58_io_data_2_in_bits),
    .io_data_2_out_valid(PE_58_io_data_2_out_valid),
    .io_data_2_out_bits(PE_58_io_data_2_out_bits),
    .io_data_1_in_valid(PE_58_io_data_1_in_valid),
    .io_data_1_in_bits(PE_58_io_data_1_in_bits),
    .io_data_1_out_valid(PE_58_io_data_1_out_valid),
    .io_data_1_out_bits(PE_58_io_data_1_out_bits),
    .io_data_0_in_valid(PE_58_io_data_0_in_valid),
    .io_data_0_in_bits(PE_58_io_data_0_in_bits),
    .io_data_0_out_valid(PE_58_io_data_0_out_valid),
    .io_data_0_out_bits(PE_58_io_data_0_out_bits),
    .io_sig_stat2trans(PE_58_io_sig_stat2trans)
  );
  PE PE_59 ( // @[pearray.scala 103:13]
    .clock(PE_59_clock),
    .reset(PE_59_reset),
    .io_data_2_in_valid(PE_59_io_data_2_in_valid),
    .io_data_2_in_bits(PE_59_io_data_2_in_bits),
    .io_data_2_out_valid(PE_59_io_data_2_out_valid),
    .io_data_2_out_bits(PE_59_io_data_2_out_bits),
    .io_data_1_in_valid(PE_59_io_data_1_in_valid),
    .io_data_1_in_bits(PE_59_io_data_1_in_bits),
    .io_data_1_out_valid(PE_59_io_data_1_out_valid),
    .io_data_1_out_bits(PE_59_io_data_1_out_bits),
    .io_data_0_in_valid(PE_59_io_data_0_in_valid),
    .io_data_0_in_bits(PE_59_io_data_0_in_bits),
    .io_data_0_out_valid(PE_59_io_data_0_out_valid),
    .io_data_0_out_bits(PE_59_io_data_0_out_bits),
    .io_sig_stat2trans(PE_59_io_sig_stat2trans)
  );
  PE PE_60 ( // @[pearray.scala 103:13]
    .clock(PE_60_clock),
    .reset(PE_60_reset),
    .io_data_2_in_valid(PE_60_io_data_2_in_valid),
    .io_data_2_in_bits(PE_60_io_data_2_in_bits),
    .io_data_2_out_valid(PE_60_io_data_2_out_valid),
    .io_data_2_out_bits(PE_60_io_data_2_out_bits),
    .io_data_1_in_valid(PE_60_io_data_1_in_valid),
    .io_data_1_in_bits(PE_60_io_data_1_in_bits),
    .io_data_1_out_valid(PE_60_io_data_1_out_valid),
    .io_data_1_out_bits(PE_60_io_data_1_out_bits),
    .io_data_0_in_valid(PE_60_io_data_0_in_valid),
    .io_data_0_in_bits(PE_60_io_data_0_in_bits),
    .io_data_0_out_valid(PE_60_io_data_0_out_valid),
    .io_data_0_out_bits(PE_60_io_data_0_out_bits),
    .io_sig_stat2trans(PE_60_io_sig_stat2trans)
  );
  PE PE_61 ( // @[pearray.scala 103:13]
    .clock(PE_61_clock),
    .reset(PE_61_reset),
    .io_data_2_in_valid(PE_61_io_data_2_in_valid),
    .io_data_2_in_bits(PE_61_io_data_2_in_bits),
    .io_data_2_out_valid(PE_61_io_data_2_out_valid),
    .io_data_2_out_bits(PE_61_io_data_2_out_bits),
    .io_data_1_in_valid(PE_61_io_data_1_in_valid),
    .io_data_1_in_bits(PE_61_io_data_1_in_bits),
    .io_data_1_out_valid(PE_61_io_data_1_out_valid),
    .io_data_1_out_bits(PE_61_io_data_1_out_bits),
    .io_data_0_in_valid(PE_61_io_data_0_in_valid),
    .io_data_0_in_bits(PE_61_io_data_0_in_bits),
    .io_data_0_out_valid(PE_61_io_data_0_out_valid),
    .io_data_0_out_bits(PE_61_io_data_0_out_bits),
    .io_sig_stat2trans(PE_61_io_sig_stat2trans)
  );
  PE PE_62 ( // @[pearray.scala 103:13]
    .clock(PE_62_clock),
    .reset(PE_62_reset),
    .io_data_2_in_valid(PE_62_io_data_2_in_valid),
    .io_data_2_in_bits(PE_62_io_data_2_in_bits),
    .io_data_2_out_valid(PE_62_io_data_2_out_valid),
    .io_data_2_out_bits(PE_62_io_data_2_out_bits),
    .io_data_1_in_valid(PE_62_io_data_1_in_valid),
    .io_data_1_in_bits(PE_62_io_data_1_in_bits),
    .io_data_1_out_valid(PE_62_io_data_1_out_valid),
    .io_data_1_out_bits(PE_62_io_data_1_out_bits),
    .io_data_0_in_valid(PE_62_io_data_0_in_valid),
    .io_data_0_in_bits(PE_62_io_data_0_in_bits),
    .io_data_0_out_valid(PE_62_io_data_0_out_valid),
    .io_data_0_out_bits(PE_62_io_data_0_out_bits),
    .io_sig_stat2trans(PE_62_io_sig_stat2trans)
  );
  PE PE_63 ( // @[pearray.scala 103:13]
    .clock(PE_63_clock),
    .reset(PE_63_reset),
    .io_data_2_in_valid(PE_63_io_data_2_in_valid),
    .io_data_2_in_bits(PE_63_io_data_2_in_bits),
    .io_data_2_out_valid(PE_63_io_data_2_out_valid),
    .io_data_2_out_bits(PE_63_io_data_2_out_bits),
    .io_data_1_in_valid(PE_63_io_data_1_in_valid),
    .io_data_1_in_bits(PE_63_io_data_1_in_bits),
    .io_data_1_out_valid(PE_63_io_data_1_out_valid),
    .io_data_1_out_bits(PE_63_io_data_1_out_bits),
    .io_data_0_in_valid(PE_63_io_data_0_in_valid),
    .io_data_0_in_bits(PE_63_io_data_0_in_bits),
    .io_data_0_out_valid(PE_63_io_data_0_out_valid),
    .io_data_0_out_bits(PE_63_io_data_0_out_bits),
    .io_sig_stat2trans(PE_63_io_sig_stat2trans)
  );
  PE PE_64 ( // @[pearray.scala 103:13]
    .clock(PE_64_clock),
    .reset(PE_64_reset),
    .io_data_2_in_valid(PE_64_io_data_2_in_valid),
    .io_data_2_in_bits(PE_64_io_data_2_in_bits),
    .io_data_2_out_valid(PE_64_io_data_2_out_valid),
    .io_data_2_out_bits(PE_64_io_data_2_out_bits),
    .io_data_1_in_valid(PE_64_io_data_1_in_valid),
    .io_data_1_in_bits(PE_64_io_data_1_in_bits),
    .io_data_1_out_valid(PE_64_io_data_1_out_valid),
    .io_data_1_out_bits(PE_64_io_data_1_out_bits),
    .io_data_0_in_valid(PE_64_io_data_0_in_valid),
    .io_data_0_in_bits(PE_64_io_data_0_in_bits),
    .io_data_0_out_valid(PE_64_io_data_0_out_valid),
    .io_data_0_out_bits(PE_64_io_data_0_out_bits),
    .io_sig_stat2trans(PE_64_io_sig_stat2trans)
  );
  PE PE_65 ( // @[pearray.scala 103:13]
    .clock(PE_65_clock),
    .reset(PE_65_reset),
    .io_data_2_in_valid(PE_65_io_data_2_in_valid),
    .io_data_2_in_bits(PE_65_io_data_2_in_bits),
    .io_data_2_out_valid(PE_65_io_data_2_out_valid),
    .io_data_2_out_bits(PE_65_io_data_2_out_bits),
    .io_data_1_in_valid(PE_65_io_data_1_in_valid),
    .io_data_1_in_bits(PE_65_io_data_1_in_bits),
    .io_data_1_out_valid(PE_65_io_data_1_out_valid),
    .io_data_1_out_bits(PE_65_io_data_1_out_bits),
    .io_data_0_in_valid(PE_65_io_data_0_in_valid),
    .io_data_0_in_bits(PE_65_io_data_0_in_bits),
    .io_data_0_out_valid(PE_65_io_data_0_out_valid),
    .io_data_0_out_bits(PE_65_io_data_0_out_bits),
    .io_sig_stat2trans(PE_65_io_sig_stat2trans)
  );
  PE PE_66 ( // @[pearray.scala 103:13]
    .clock(PE_66_clock),
    .reset(PE_66_reset),
    .io_data_2_in_valid(PE_66_io_data_2_in_valid),
    .io_data_2_in_bits(PE_66_io_data_2_in_bits),
    .io_data_2_out_valid(PE_66_io_data_2_out_valid),
    .io_data_2_out_bits(PE_66_io_data_2_out_bits),
    .io_data_1_in_valid(PE_66_io_data_1_in_valid),
    .io_data_1_in_bits(PE_66_io_data_1_in_bits),
    .io_data_1_out_valid(PE_66_io_data_1_out_valid),
    .io_data_1_out_bits(PE_66_io_data_1_out_bits),
    .io_data_0_in_valid(PE_66_io_data_0_in_valid),
    .io_data_0_in_bits(PE_66_io_data_0_in_bits),
    .io_data_0_out_valid(PE_66_io_data_0_out_valid),
    .io_data_0_out_bits(PE_66_io_data_0_out_bits),
    .io_sig_stat2trans(PE_66_io_sig_stat2trans)
  );
  PE PE_67 ( // @[pearray.scala 103:13]
    .clock(PE_67_clock),
    .reset(PE_67_reset),
    .io_data_2_in_valid(PE_67_io_data_2_in_valid),
    .io_data_2_in_bits(PE_67_io_data_2_in_bits),
    .io_data_2_out_valid(PE_67_io_data_2_out_valid),
    .io_data_2_out_bits(PE_67_io_data_2_out_bits),
    .io_data_1_in_valid(PE_67_io_data_1_in_valid),
    .io_data_1_in_bits(PE_67_io_data_1_in_bits),
    .io_data_1_out_valid(PE_67_io_data_1_out_valid),
    .io_data_1_out_bits(PE_67_io_data_1_out_bits),
    .io_data_0_in_valid(PE_67_io_data_0_in_valid),
    .io_data_0_in_bits(PE_67_io_data_0_in_bits),
    .io_data_0_out_valid(PE_67_io_data_0_out_valid),
    .io_data_0_out_bits(PE_67_io_data_0_out_bits),
    .io_sig_stat2trans(PE_67_io_sig_stat2trans)
  );
  PE PE_68 ( // @[pearray.scala 103:13]
    .clock(PE_68_clock),
    .reset(PE_68_reset),
    .io_data_2_in_valid(PE_68_io_data_2_in_valid),
    .io_data_2_in_bits(PE_68_io_data_2_in_bits),
    .io_data_2_out_valid(PE_68_io_data_2_out_valid),
    .io_data_2_out_bits(PE_68_io_data_2_out_bits),
    .io_data_1_in_valid(PE_68_io_data_1_in_valid),
    .io_data_1_in_bits(PE_68_io_data_1_in_bits),
    .io_data_1_out_valid(PE_68_io_data_1_out_valid),
    .io_data_1_out_bits(PE_68_io_data_1_out_bits),
    .io_data_0_in_valid(PE_68_io_data_0_in_valid),
    .io_data_0_in_bits(PE_68_io_data_0_in_bits),
    .io_data_0_out_valid(PE_68_io_data_0_out_valid),
    .io_data_0_out_bits(PE_68_io_data_0_out_bits),
    .io_sig_stat2trans(PE_68_io_sig_stat2trans)
  );
  PE PE_69 ( // @[pearray.scala 103:13]
    .clock(PE_69_clock),
    .reset(PE_69_reset),
    .io_data_2_in_valid(PE_69_io_data_2_in_valid),
    .io_data_2_in_bits(PE_69_io_data_2_in_bits),
    .io_data_2_out_valid(PE_69_io_data_2_out_valid),
    .io_data_2_out_bits(PE_69_io_data_2_out_bits),
    .io_data_1_in_valid(PE_69_io_data_1_in_valid),
    .io_data_1_in_bits(PE_69_io_data_1_in_bits),
    .io_data_1_out_valid(PE_69_io_data_1_out_valid),
    .io_data_1_out_bits(PE_69_io_data_1_out_bits),
    .io_data_0_in_valid(PE_69_io_data_0_in_valid),
    .io_data_0_in_bits(PE_69_io_data_0_in_bits),
    .io_data_0_out_valid(PE_69_io_data_0_out_valid),
    .io_data_0_out_bits(PE_69_io_data_0_out_bits),
    .io_sig_stat2trans(PE_69_io_sig_stat2trans)
  );
  PE PE_70 ( // @[pearray.scala 103:13]
    .clock(PE_70_clock),
    .reset(PE_70_reset),
    .io_data_2_in_valid(PE_70_io_data_2_in_valid),
    .io_data_2_in_bits(PE_70_io_data_2_in_bits),
    .io_data_2_out_valid(PE_70_io_data_2_out_valid),
    .io_data_2_out_bits(PE_70_io_data_2_out_bits),
    .io_data_1_in_valid(PE_70_io_data_1_in_valid),
    .io_data_1_in_bits(PE_70_io_data_1_in_bits),
    .io_data_1_out_valid(PE_70_io_data_1_out_valid),
    .io_data_1_out_bits(PE_70_io_data_1_out_bits),
    .io_data_0_in_valid(PE_70_io_data_0_in_valid),
    .io_data_0_in_bits(PE_70_io_data_0_in_bits),
    .io_data_0_out_valid(PE_70_io_data_0_out_valid),
    .io_data_0_out_bits(PE_70_io_data_0_out_bits),
    .io_sig_stat2trans(PE_70_io_sig_stat2trans)
  );
  PE PE_71 ( // @[pearray.scala 103:13]
    .clock(PE_71_clock),
    .reset(PE_71_reset),
    .io_data_2_in_valid(PE_71_io_data_2_in_valid),
    .io_data_2_in_bits(PE_71_io_data_2_in_bits),
    .io_data_2_out_valid(PE_71_io_data_2_out_valid),
    .io_data_2_out_bits(PE_71_io_data_2_out_bits),
    .io_data_1_in_valid(PE_71_io_data_1_in_valid),
    .io_data_1_in_bits(PE_71_io_data_1_in_bits),
    .io_data_1_out_valid(PE_71_io_data_1_out_valid),
    .io_data_1_out_bits(PE_71_io_data_1_out_bits),
    .io_data_0_in_valid(PE_71_io_data_0_in_valid),
    .io_data_0_in_bits(PE_71_io_data_0_in_bits),
    .io_data_0_out_valid(PE_71_io_data_0_out_valid),
    .io_data_0_out_bits(PE_71_io_data_0_out_bits),
    .io_sig_stat2trans(PE_71_io_sig_stat2trans)
  );
  PE PE_72 ( // @[pearray.scala 103:13]
    .clock(PE_72_clock),
    .reset(PE_72_reset),
    .io_data_2_in_valid(PE_72_io_data_2_in_valid),
    .io_data_2_in_bits(PE_72_io_data_2_in_bits),
    .io_data_2_out_valid(PE_72_io_data_2_out_valid),
    .io_data_2_out_bits(PE_72_io_data_2_out_bits),
    .io_data_1_in_valid(PE_72_io_data_1_in_valid),
    .io_data_1_in_bits(PE_72_io_data_1_in_bits),
    .io_data_1_out_valid(PE_72_io_data_1_out_valid),
    .io_data_1_out_bits(PE_72_io_data_1_out_bits),
    .io_data_0_in_valid(PE_72_io_data_0_in_valid),
    .io_data_0_in_bits(PE_72_io_data_0_in_bits),
    .io_data_0_out_valid(PE_72_io_data_0_out_valid),
    .io_data_0_out_bits(PE_72_io_data_0_out_bits),
    .io_sig_stat2trans(PE_72_io_sig_stat2trans)
  );
  PE PE_73 ( // @[pearray.scala 103:13]
    .clock(PE_73_clock),
    .reset(PE_73_reset),
    .io_data_2_in_valid(PE_73_io_data_2_in_valid),
    .io_data_2_in_bits(PE_73_io_data_2_in_bits),
    .io_data_2_out_valid(PE_73_io_data_2_out_valid),
    .io_data_2_out_bits(PE_73_io_data_2_out_bits),
    .io_data_1_in_valid(PE_73_io_data_1_in_valid),
    .io_data_1_in_bits(PE_73_io_data_1_in_bits),
    .io_data_1_out_valid(PE_73_io_data_1_out_valid),
    .io_data_1_out_bits(PE_73_io_data_1_out_bits),
    .io_data_0_in_valid(PE_73_io_data_0_in_valid),
    .io_data_0_in_bits(PE_73_io_data_0_in_bits),
    .io_data_0_out_valid(PE_73_io_data_0_out_valid),
    .io_data_0_out_bits(PE_73_io_data_0_out_bits),
    .io_sig_stat2trans(PE_73_io_sig_stat2trans)
  );
  PE PE_74 ( // @[pearray.scala 103:13]
    .clock(PE_74_clock),
    .reset(PE_74_reset),
    .io_data_2_in_valid(PE_74_io_data_2_in_valid),
    .io_data_2_in_bits(PE_74_io_data_2_in_bits),
    .io_data_2_out_valid(PE_74_io_data_2_out_valid),
    .io_data_2_out_bits(PE_74_io_data_2_out_bits),
    .io_data_1_in_valid(PE_74_io_data_1_in_valid),
    .io_data_1_in_bits(PE_74_io_data_1_in_bits),
    .io_data_1_out_valid(PE_74_io_data_1_out_valid),
    .io_data_1_out_bits(PE_74_io_data_1_out_bits),
    .io_data_0_in_valid(PE_74_io_data_0_in_valid),
    .io_data_0_in_bits(PE_74_io_data_0_in_bits),
    .io_data_0_out_valid(PE_74_io_data_0_out_valid),
    .io_data_0_out_bits(PE_74_io_data_0_out_bits),
    .io_sig_stat2trans(PE_74_io_sig_stat2trans)
  );
  PE PE_75 ( // @[pearray.scala 103:13]
    .clock(PE_75_clock),
    .reset(PE_75_reset),
    .io_data_2_in_valid(PE_75_io_data_2_in_valid),
    .io_data_2_in_bits(PE_75_io_data_2_in_bits),
    .io_data_2_out_valid(PE_75_io_data_2_out_valid),
    .io_data_2_out_bits(PE_75_io_data_2_out_bits),
    .io_data_1_in_valid(PE_75_io_data_1_in_valid),
    .io_data_1_in_bits(PE_75_io_data_1_in_bits),
    .io_data_1_out_valid(PE_75_io_data_1_out_valid),
    .io_data_1_out_bits(PE_75_io_data_1_out_bits),
    .io_data_0_in_valid(PE_75_io_data_0_in_valid),
    .io_data_0_in_bits(PE_75_io_data_0_in_bits),
    .io_data_0_out_valid(PE_75_io_data_0_out_valid),
    .io_data_0_out_bits(PE_75_io_data_0_out_bits),
    .io_sig_stat2trans(PE_75_io_sig_stat2trans)
  );
  PE PE_76 ( // @[pearray.scala 103:13]
    .clock(PE_76_clock),
    .reset(PE_76_reset),
    .io_data_2_in_valid(PE_76_io_data_2_in_valid),
    .io_data_2_in_bits(PE_76_io_data_2_in_bits),
    .io_data_2_out_valid(PE_76_io_data_2_out_valid),
    .io_data_2_out_bits(PE_76_io_data_2_out_bits),
    .io_data_1_in_valid(PE_76_io_data_1_in_valid),
    .io_data_1_in_bits(PE_76_io_data_1_in_bits),
    .io_data_1_out_valid(PE_76_io_data_1_out_valid),
    .io_data_1_out_bits(PE_76_io_data_1_out_bits),
    .io_data_0_in_valid(PE_76_io_data_0_in_valid),
    .io_data_0_in_bits(PE_76_io_data_0_in_bits),
    .io_data_0_out_valid(PE_76_io_data_0_out_valid),
    .io_data_0_out_bits(PE_76_io_data_0_out_bits),
    .io_sig_stat2trans(PE_76_io_sig_stat2trans)
  );
  PE PE_77 ( // @[pearray.scala 103:13]
    .clock(PE_77_clock),
    .reset(PE_77_reset),
    .io_data_2_in_valid(PE_77_io_data_2_in_valid),
    .io_data_2_in_bits(PE_77_io_data_2_in_bits),
    .io_data_2_out_valid(PE_77_io_data_2_out_valid),
    .io_data_2_out_bits(PE_77_io_data_2_out_bits),
    .io_data_1_in_valid(PE_77_io_data_1_in_valid),
    .io_data_1_in_bits(PE_77_io_data_1_in_bits),
    .io_data_1_out_valid(PE_77_io_data_1_out_valid),
    .io_data_1_out_bits(PE_77_io_data_1_out_bits),
    .io_data_0_in_valid(PE_77_io_data_0_in_valid),
    .io_data_0_in_bits(PE_77_io_data_0_in_bits),
    .io_data_0_out_valid(PE_77_io_data_0_out_valid),
    .io_data_0_out_bits(PE_77_io_data_0_out_bits),
    .io_sig_stat2trans(PE_77_io_sig_stat2trans)
  );
  PE PE_78 ( // @[pearray.scala 103:13]
    .clock(PE_78_clock),
    .reset(PE_78_reset),
    .io_data_2_in_valid(PE_78_io_data_2_in_valid),
    .io_data_2_in_bits(PE_78_io_data_2_in_bits),
    .io_data_2_out_valid(PE_78_io_data_2_out_valid),
    .io_data_2_out_bits(PE_78_io_data_2_out_bits),
    .io_data_1_in_valid(PE_78_io_data_1_in_valid),
    .io_data_1_in_bits(PE_78_io_data_1_in_bits),
    .io_data_1_out_valid(PE_78_io_data_1_out_valid),
    .io_data_1_out_bits(PE_78_io_data_1_out_bits),
    .io_data_0_in_valid(PE_78_io_data_0_in_valid),
    .io_data_0_in_bits(PE_78_io_data_0_in_bits),
    .io_data_0_out_valid(PE_78_io_data_0_out_valid),
    .io_data_0_out_bits(PE_78_io_data_0_out_bits),
    .io_sig_stat2trans(PE_78_io_sig_stat2trans)
  );
  PE PE_79 ( // @[pearray.scala 103:13]
    .clock(PE_79_clock),
    .reset(PE_79_reset),
    .io_data_2_in_valid(PE_79_io_data_2_in_valid),
    .io_data_2_in_bits(PE_79_io_data_2_in_bits),
    .io_data_2_out_valid(PE_79_io_data_2_out_valid),
    .io_data_2_out_bits(PE_79_io_data_2_out_bits),
    .io_data_1_in_valid(PE_79_io_data_1_in_valid),
    .io_data_1_in_bits(PE_79_io_data_1_in_bits),
    .io_data_1_out_valid(PE_79_io_data_1_out_valid),
    .io_data_1_out_bits(PE_79_io_data_1_out_bits),
    .io_data_0_in_valid(PE_79_io_data_0_in_valid),
    .io_data_0_in_bits(PE_79_io_data_0_in_bits),
    .io_data_0_out_valid(PE_79_io_data_0_out_valid),
    .io_data_0_out_bits(PE_79_io_data_0_out_bits),
    .io_sig_stat2trans(PE_79_io_sig_stat2trans)
  );
  PE PE_80 ( // @[pearray.scala 103:13]
    .clock(PE_80_clock),
    .reset(PE_80_reset),
    .io_data_2_in_valid(PE_80_io_data_2_in_valid),
    .io_data_2_in_bits(PE_80_io_data_2_in_bits),
    .io_data_2_out_valid(PE_80_io_data_2_out_valid),
    .io_data_2_out_bits(PE_80_io_data_2_out_bits),
    .io_data_1_in_valid(PE_80_io_data_1_in_valid),
    .io_data_1_in_bits(PE_80_io_data_1_in_bits),
    .io_data_1_out_valid(PE_80_io_data_1_out_valid),
    .io_data_1_out_bits(PE_80_io_data_1_out_bits),
    .io_data_0_in_valid(PE_80_io_data_0_in_valid),
    .io_data_0_in_bits(PE_80_io_data_0_in_bits),
    .io_data_0_out_valid(PE_80_io_data_0_out_valid),
    .io_data_0_out_bits(PE_80_io_data_0_out_bits),
    .io_sig_stat2trans(PE_80_io_sig_stat2trans)
  );
  PE PE_81 ( // @[pearray.scala 103:13]
    .clock(PE_81_clock),
    .reset(PE_81_reset),
    .io_data_2_in_valid(PE_81_io_data_2_in_valid),
    .io_data_2_in_bits(PE_81_io_data_2_in_bits),
    .io_data_2_out_valid(PE_81_io_data_2_out_valid),
    .io_data_2_out_bits(PE_81_io_data_2_out_bits),
    .io_data_1_in_valid(PE_81_io_data_1_in_valid),
    .io_data_1_in_bits(PE_81_io_data_1_in_bits),
    .io_data_1_out_valid(PE_81_io_data_1_out_valid),
    .io_data_1_out_bits(PE_81_io_data_1_out_bits),
    .io_data_0_in_valid(PE_81_io_data_0_in_valid),
    .io_data_0_in_bits(PE_81_io_data_0_in_bits),
    .io_data_0_out_valid(PE_81_io_data_0_out_valid),
    .io_data_0_out_bits(PE_81_io_data_0_out_bits),
    .io_sig_stat2trans(PE_81_io_sig_stat2trans)
  );
  PE PE_82 ( // @[pearray.scala 103:13]
    .clock(PE_82_clock),
    .reset(PE_82_reset),
    .io_data_2_in_valid(PE_82_io_data_2_in_valid),
    .io_data_2_in_bits(PE_82_io_data_2_in_bits),
    .io_data_2_out_valid(PE_82_io_data_2_out_valid),
    .io_data_2_out_bits(PE_82_io_data_2_out_bits),
    .io_data_1_in_valid(PE_82_io_data_1_in_valid),
    .io_data_1_in_bits(PE_82_io_data_1_in_bits),
    .io_data_1_out_valid(PE_82_io_data_1_out_valid),
    .io_data_1_out_bits(PE_82_io_data_1_out_bits),
    .io_data_0_in_valid(PE_82_io_data_0_in_valid),
    .io_data_0_in_bits(PE_82_io_data_0_in_bits),
    .io_data_0_out_valid(PE_82_io_data_0_out_valid),
    .io_data_0_out_bits(PE_82_io_data_0_out_bits),
    .io_sig_stat2trans(PE_82_io_sig_stat2trans)
  );
  PE PE_83 ( // @[pearray.scala 103:13]
    .clock(PE_83_clock),
    .reset(PE_83_reset),
    .io_data_2_in_valid(PE_83_io_data_2_in_valid),
    .io_data_2_in_bits(PE_83_io_data_2_in_bits),
    .io_data_2_out_valid(PE_83_io_data_2_out_valid),
    .io_data_2_out_bits(PE_83_io_data_2_out_bits),
    .io_data_1_in_valid(PE_83_io_data_1_in_valid),
    .io_data_1_in_bits(PE_83_io_data_1_in_bits),
    .io_data_1_out_valid(PE_83_io_data_1_out_valid),
    .io_data_1_out_bits(PE_83_io_data_1_out_bits),
    .io_data_0_in_valid(PE_83_io_data_0_in_valid),
    .io_data_0_in_bits(PE_83_io_data_0_in_bits),
    .io_data_0_out_valid(PE_83_io_data_0_out_valid),
    .io_data_0_out_bits(PE_83_io_data_0_out_bits),
    .io_sig_stat2trans(PE_83_io_sig_stat2trans)
  );
  PE PE_84 ( // @[pearray.scala 103:13]
    .clock(PE_84_clock),
    .reset(PE_84_reset),
    .io_data_2_in_valid(PE_84_io_data_2_in_valid),
    .io_data_2_in_bits(PE_84_io_data_2_in_bits),
    .io_data_2_out_valid(PE_84_io_data_2_out_valid),
    .io_data_2_out_bits(PE_84_io_data_2_out_bits),
    .io_data_1_in_valid(PE_84_io_data_1_in_valid),
    .io_data_1_in_bits(PE_84_io_data_1_in_bits),
    .io_data_1_out_valid(PE_84_io_data_1_out_valid),
    .io_data_1_out_bits(PE_84_io_data_1_out_bits),
    .io_data_0_in_valid(PE_84_io_data_0_in_valid),
    .io_data_0_in_bits(PE_84_io_data_0_in_bits),
    .io_data_0_out_valid(PE_84_io_data_0_out_valid),
    .io_data_0_out_bits(PE_84_io_data_0_out_bits),
    .io_sig_stat2trans(PE_84_io_sig_stat2trans)
  );
  PE PE_85 ( // @[pearray.scala 103:13]
    .clock(PE_85_clock),
    .reset(PE_85_reset),
    .io_data_2_in_valid(PE_85_io_data_2_in_valid),
    .io_data_2_in_bits(PE_85_io_data_2_in_bits),
    .io_data_2_out_valid(PE_85_io_data_2_out_valid),
    .io_data_2_out_bits(PE_85_io_data_2_out_bits),
    .io_data_1_in_valid(PE_85_io_data_1_in_valid),
    .io_data_1_in_bits(PE_85_io_data_1_in_bits),
    .io_data_1_out_valid(PE_85_io_data_1_out_valid),
    .io_data_1_out_bits(PE_85_io_data_1_out_bits),
    .io_data_0_in_valid(PE_85_io_data_0_in_valid),
    .io_data_0_in_bits(PE_85_io_data_0_in_bits),
    .io_data_0_out_valid(PE_85_io_data_0_out_valid),
    .io_data_0_out_bits(PE_85_io_data_0_out_bits),
    .io_sig_stat2trans(PE_85_io_sig_stat2trans)
  );
  PE PE_86 ( // @[pearray.scala 103:13]
    .clock(PE_86_clock),
    .reset(PE_86_reset),
    .io_data_2_in_valid(PE_86_io_data_2_in_valid),
    .io_data_2_in_bits(PE_86_io_data_2_in_bits),
    .io_data_2_out_valid(PE_86_io_data_2_out_valid),
    .io_data_2_out_bits(PE_86_io_data_2_out_bits),
    .io_data_1_in_valid(PE_86_io_data_1_in_valid),
    .io_data_1_in_bits(PE_86_io_data_1_in_bits),
    .io_data_1_out_valid(PE_86_io_data_1_out_valid),
    .io_data_1_out_bits(PE_86_io_data_1_out_bits),
    .io_data_0_in_valid(PE_86_io_data_0_in_valid),
    .io_data_0_in_bits(PE_86_io_data_0_in_bits),
    .io_data_0_out_valid(PE_86_io_data_0_out_valid),
    .io_data_0_out_bits(PE_86_io_data_0_out_bits),
    .io_sig_stat2trans(PE_86_io_sig_stat2trans)
  );
  PE PE_87 ( // @[pearray.scala 103:13]
    .clock(PE_87_clock),
    .reset(PE_87_reset),
    .io_data_2_in_valid(PE_87_io_data_2_in_valid),
    .io_data_2_in_bits(PE_87_io_data_2_in_bits),
    .io_data_2_out_valid(PE_87_io_data_2_out_valid),
    .io_data_2_out_bits(PE_87_io_data_2_out_bits),
    .io_data_1_in_valid(PE_87_io_data_1_in_valid),
    .io_data_1_in_bits(PE_87_io_data_1_in_bits),
    .io_data_1_out_valid(PE_87_io_data_1_out_valid),
    .io_data_1_out_bits(PE_87_io_data_1_out_bits),
    .io_data_0_in_valid(PE_87_io_data_0_in_valid),
    .io_data_0_in_bits(PE_87_io_data_0_in_bits),
    .io_data_0_out_valid(PE_87_io_data_0_out_valid),
    .io_data_0_out_bits(PE_87_io_data_0_out_bits),
    .io_sig_stat2trans(PE_87_io_sig_stat2trans)
  );
  PE PE_88 ( // @[pearray.scala 103:13]
    .clock(PE_88_clock),
    .reset(PE_88_reset),
    .io_data_2_in_valid(PE_88_io_data_2_in_valid),
    .io_data_2_in_bits(PE_88_io_data_2_in_bits),
    .io_data_2_out_valid(PE_88_io_data_2_out_valid),
    .io_data_2_out_bits(PE_88_io_data_2_out_bits),
    .io_data_1_in_valid(PE_88_io_data_1_in_valid),
    .io_data_1_in_bits(PE_88_io_data_1_in_bits),
    .io_data_1_out_valid(PE_88_io_data_1_out_valid),
    .io_data_1_out_bits(PE_88_io_data_1_out_bits),
    .io_data_0_in_valid(PE_88_io_data_0_in_valid),
    .io_data_0_in_bits(PE_88_io_data_0_in_bits),
    .io_data_0_out_valid(PE_88_io_data_0_out_valid),
    .io_data_0_out_bits(PE_88_io_data_0_out_bits),
    .io_sig_stat2trans(PE_88_io_sig_stat2trans)
  );
  PE PE_89 ( // @[pearray.scala 103:13]
    .clock(PE_89_clock),
    .reset(PE_89_reset),
    .io_data_2_in_valid(PE_89_io_data_2_in_valid),
    .io_data_2_in_bits(PE_89_io_data_2_in_bits),
    .io_data_2_out_valid(PE_89_io_data_2_out_valid),
    .io_data_2_out_bits(PE_89_io_data_2_out_bits),
    .io_data_1_in_valid(PE_89_io_data_1_in_valid),
    .io_data_1_in_bits(PE_89_io_data_1_in_bits),
    .io_data_1_out_valid(PE_89_io_data_1_out_valid),
    .io_data_1_out_bits(PE_89_io_data_1_out_bits),
    .io_data_0_in_valid(PE_89_io_data_0_in_valid),
    .io_data_0_in_bits(PE_89_io_data_0_in_bits),
    .io_data_0_out_valid(PE_89_io_data_0_out_valid),
    .io_data_0_out_bits(PE_89_io_data_0_out_bits),
    .io_sig_stat2trans(PE_89_io_sig_stat2trans)
  );
  PE PE_90 ( // @[pearray.scala 103:13]
    .clock(PE_90_clock),
    .reset(PE_90_reset),
    .io_data_2_in_valid(PE_90_io_data_2_in_valid),
    .io_data_2_in_bits(PE_90_io_data_2_in_bits),
    .io_data_2_out_valid(PE_90_io_data_2_out_valid),
    .io_data_2_out_bits(PE_90_io_data_2_out_bits),
    .io_data_1_in_valid(PE_90_io_data_1_in_valid),
    .io_data_1_in_bits(PE_90_io_data_1_in_bits),
    .io_data_1_out_valid(PE_90_io_data_1_out_valid),
    .io_data_1_out_bits(PE_90_io_data_1_out_bits),
    .io_data_0_in_valid(PE_90_io_data_0_in_valid),
    .io_data_0_in_bits(PE_90_io_data_0_in_bits),
    .io_data_0_out_valid(PE_90_io_data_0_out_valid),
    .io_data_0_out_bits(PE_90_io_data_0_out_bits),
    .io_sig_stat2trans(PE_90_io_sig_stat2trans)
  );
  PE PE_91 ( // @[pearray.scala 103:13]
    .clock(PE_91_clock),
    .reset(PE_91_reset),
    .io_data_2_in_valid(PE_91_io_data_2_in_valid),
    .io_data_2_in_bits(PE_91_io_data_2_in_bits),
    .io_data_2_out_valid(PE_91_io_data_2_out_valid),
    .io_data_2_out_bits(PE_91_io_data_2_out_bits),
    .io_data_1_in_valid(PE_91_io_data_1_in_valid),
    .io_data_1_in_bits(PE_91_io_data_1_in_bits),
    .io_data_1_out_valid(PE_91_io_data_1_out_valid),
    .io_data_1_out_bits(PE_91_io_data_1_out_bits),
    .io_data_0_in_valid(PE_91_io_data_0_in_valid),
    .io_data_0_in_bits(PE_91_io_data_0_in_bits),
    .io_data_0_out_valid(PE_91_io_data_0_out_valid),
    .io_data_0_out_bits(PE_91_io_data_0_out_bits),
    .io_sig_stat2trans(PE_91_io_sig_stat2trans)
  );
  PE PE_92 ( // @[pearray.scala 103:13]
    .clock(PE_92_clock),
    .reset(PE_92_reset),
    .io_data_2_in_valid(PE_92_io_data_2_in_valid),
    .io_data_2_in_bits(PE_92_io_data_2_in_bits),
    .io_data_2_out_valid(PE_92_io_data_2_out_valid),
    .io_data_2_out_bits(PE_92_io_data_2_out_bits),
    .io_data_1_in_valid(PE_92_io_data_1_in_valid),
    .io_data_1_in_bits(PE_92_io_data_1_in_bits),
    .io_data_1_out_valid(PE_92_io_data_1_out_valid),
    .io_data_1_out_bits(PE_92_io_data_1_out_bits),
    .io_data_0_in_valid(PE_92_io_data_0_in_valid),
    .io_data_0_in_bits(PE_92_io_data_0_in_bits),
    .io_data_0_out_valid(PE_92_io_data_0_out_valid),
    .io_data_0_out_bits(PE_92_io_data_0_out_bits),
    .io_sig_stat2trans(PE_92_io_sig_stat2trans)
  );
  PE PE_93 ( // @[pearray.scala 103:13]
    .clock(PE_93_clock),
    .reset(PE_93_reset),
    .io_data_2_in_valid(PE_93_io_data_2_in_valid),
    .io_data_2_in_bits(PE_93_io_data_2_in_bits),
    .io_data_2_out_valid(PE_93_io_data_2_out_valid),
    .io_data_2_out_bits(PE_93_io_data_2_out_bits),
    .io_data_1_in_valid(PE_93_io_data_1_in_valid),
    .io_data_1_in_bits(PE_93_io_data_1_in_bits),
    .io_data_1_out_valid(PE_93_io_data_1_out_valid),
    .io_data_1_out_bits(PE_93_io_data_1_out_bits),
    .io_data_0_in_valid(PE_93_io_data_0_in_valid),
    .io_data_0_in_bits(PE_93_io_data_0_in_bits),
    .io_data_0_out_valid(PE_93_io_data_0_out_valid),
    .io_data_0_out_bits(PE_93_io_data_0_out_bits),
    .io_sig_stat2trans(PE_93_io_sig_stat2trans)
  );
  PE PE_94 ( // @[pearray.scala 103:13]
    .clock(PE_94_clock),
    .reset(PE_94_reset),
    .io_data_2_in_valid(PE_94_io_data_2_in_valid),
    .io_data_2_in_bits(PE_94_io_data_2_in_bits),
    .io_data_2_out_valid(PE_94_io_data_2_out_valid),
    .io_data_2_out_bits(PE_94_io_data_2_out_bits),
    .io_data_1_in_valid(PE_94_io_data_1_in_valid),
    .io_data_1_in_bits(PE_94_io_data_1_in_bits),
    .io_data_1_out_valid(PE_94_io_data_1_out_valid),
    .io_data_1_out_bits(PE_94_io_data_1_out_bits),
    .io_data_0_in_valid(PE_94_io_data_0_in_valid),
    .io_data_0_in_bits(PE_94_io_data_0_in_bits),
    .io_data_0_out_valid(PE_94_io_data_0_out_valid),
    .io_data_0_out_bits(PE_94_io_data_0_out_bits),
    .io_sig_stat2trans(PE_94_io_sig_stat2trans)
  );
  PE PE_95 ( // @[pearray.scala 103:13]
    .clock(PE_95_clock),
    .reset(PE_95_reset),
    .io_data_2_in_valid(PE_95_io_data_2_in_valid),
    .io_data_2_in_bits(PE_95_io_data_2_in_bits),
    .io_data_2_out_valid(PE_95_io_data_2_out_valid),
    .io_data_2_out_bits(PE_95_io_data_2_out_bits),
    .io_data_1_in_valid(PE_95_io_data_1_in_valid),
    .io_data_1_in_bits(PE_95_io_data_1_in_bits),
    .io_data_1_out_valid(PE_95_io_data_1_out_valid),
    .io_data_1_out_bits(PE_95_io_data_1_out_bits),
    .io_data_0_in_valid(PE_95_io_data_0_in_valid),
    .io_data_0_in_bits(PE_95_io_data_0_in_bits),
    .io_data_0_out_valid(PE_95_io_data_0_out_valid),
    .io_data_0_out_bits(PE_95_io_data_0_out_bits),
    .io_sig_stat2trans(PE_95_io_sig_stat2trans)
  );
  PE PE_96 ( // @[pearray.scala 103:13]
    .clock(PE_96_clock),
    .reset(PE_96_reset),
    .io_data_2_in_valid(PE_96_io_data_2_in_valid),
    .io_data_2_in_bits(PE_96_io_data_2_in_bits),
    .io_data_2_out_valid(PE_96_io_data_2_out_valid),
    .io_data_2_out_bits(PE_96_io_data_2_out_bits),
    .io_data_1_in_valid(PE_96_io_data_1_in_valid),
    .io_data_1_in_bits(PE_96_io_data_1_in_bits),
    .io_data_1_out_valid(PE_96_io_data_1_out_valid),
    .io_data_1_out_bits(PE_96_io_data_1_out_bits),
    .io_data_0_in_valid(PE_96_io_data_0_in_valid),
    .io_data_0_in_bits(PE_96_io_data_0_in_bits),
    .io_data_0_out_valid(PE_96_io_data_0_out_valid),
    .io_data_0_out_bits(PE_96_io_data_0_out_bits),
    .io_sig_stat2trans(PE_96_io_sig_stat2trans)
  );
  PE PE_97 ( // @[pearray.scala 103:13]
    .clock(PE_97_clock),
    .reset(PE_97_reset),
    .io_data_2_in_valid(PE_97_io_data_2_in_valid),
    .io_data_2_in_bits(PE_97_io_data_2_in_bits),
    .io_data_2_out_valid(PE_97_io_data_2_out_valid),
    .io_data_2_out_bits(PE_97_io_data_2_out_bits),
    .io_data_1_in_valid(PE_97_io_data_1_in_valid),
    .io_data_1_in_bits(PE_97_io_data_1_in_bits),
    .io_data_1_out_valid(PE_97_io_data_1_out_valid),
    .io_data_1_out_bits(PE_97_io_data_1_out_bits),
    .io_data_0_in_valid(PE_97_io_data_0_in_valid),
    .io_data_0_in_bits(PE_97_io_data_0_in_bits),
    .io_data_0_out_valid(PE_97_io_data_0_out_valid),
    .io_data_0_out_bits(PE_97_io_data_0_out_bits),
    .io_sig_stat2trans(PE_97_io_sig_stat2trans)
  );
  PE PE_98 ( // @[pearray.scala 103:13]
    .clock(PE_98_clock),
    .reset(PE_98_reset),
    .io_data_2_in_valid(PE_98_io_data_2_in_valid),
    .io_data_2_in_bits(PE_98_io_data_2_in_bits),
    .io_data_2_out_valid(PE_98_io_data_2_out_valid),
    .io_data_2_out_bits(PE_98_io_data_2_out_bits),
    .io_data_1_in_valid(PE_98_io_data_1_in_valid),
    .io_data_1_in_bits(PE_98_io_data_1_in_bits),
    .io_data_1_out_valid(PE_98_io_data_1_out_valid),
    .io_data_1_out_bits(PE_98_io_data_1_out_bits),
    .io_data_0_in_valid(PE_98_io_data_0_in_valid),
    .io_data_0_in_bits(PE_98_io_data_0_in_bits),
    .io_data_0_out_valid(PE_98_io_data_0_out_valid),
    .io_data_0_out_bits(PE_98_io_data_0_out_bits),
    .io_sig_stat2trans(PE_98_io_sig_stat2trans)
  );
  PE PE_99 ( // @[pearray.scala 103:13]
    .clock(PE_99_clock),
    .reset(PE_99_reset),
    .io_data_2_in_valid(PE_99_io_data_2_in_valid),
    .io_data_2_in_bits(PE_99_io_data_2_in_bits),
    .io_data_2_out_valid(PE_99_io_data_2_out_valid),
    .io_data_2_out_bits(PE_99_io_data_2_out_bits),
    .io_data_1_in_valid(PE_99_io_data_1_in_valid),
    .io_data_1_in_bits(PE_99_io_data_1_in_bits),
    .io_data_1_out_valid(PE_99_io_data_1_out_valid),
    .io_data_1_out_bits(PE_99_io_data_1_out_bits),
    .io_data_0_in_valid(PE_99_io_data_0_in_valid),
    .io_data_0_in_bits(PE_99_io_data_0_in_bits),
    .io_data_0_out_valid(PE_99_io_data_0_out_valid),
    .io_data_0_out_bits(PE_99_io_data_0_out_bits),
    .io_sig_stat2trans(PE_99_io_sig_stat2trans)
  );
  PE PE_100 ( // @[pearray.scala 103:13]
    .clock(PE_100_clock),
    .reset(PE_100_reset),
    .io_data_2_in_valid(PE_100_io_data_2_in_valid),
    .io_data_2_in_bits(PE_100_io_data_2_in_bits),
    .io_data_2_out_valid(PE_100_io_data_2_out_valid),
    .io_data_2_out_bits(PE_100_io_data_2_out_bits),
    .io_data_1_in_valid(PE_100_io_data_1_in_valid),
    .io_data_1_in_bits(PE_100_io_data_1_in_bits),
    .io_data_1_out_valid(PE_100_io_data_1_out_valid),
    .io_data_1_out_bits(PE_100_io_data_1_out_bits),
    .io_data_0_in_valid(PE_100_io_data_0_in_valid),
    .io_data_0_in_bits(PE_100_io_data_0_in_bits),
    .io_data_0_out_valid(PE_100_io_data_0_out_valid),
    .io_data_0_out_bits(PE_100_io_data_0_out_bits),
    .io_sig_stat2trans(PE_100_io_sig_stat2trans)
  );
  PE PE_101 ( // @[pearray.scala 103:13]
    .clock(PE_101_clock),
    .reset(PE_101_reset),
    .io_data_2_in_valid(PE_101_io_data_2_in_valid),
    .io_data_2_in_bits(PE_101_io_data_2_in_bits),
    .io_data_2_out_valid(PE_101_io_data_2_out_valid),
    .io_data_2_out_bits(PE_101_io_data_2_out_bits),
    .io_data_1_in_valid(PE_101_io_data_1_in_valid),
    .io_data_1_in_bits(PE_101_io_data_1_in_bits),
    .io_data_1_out_valid(PE_101_io_data_1_out_valid),
    .io_data_1_out_bits(PE_101_io_data_1_out_bits),
    .io_data_0_in_valid(PE_101_io_data_0_in_valid),
    .io_data_0_in_bits(PE_101_io_data_0_in_bits),
    .io_data_0_out_valid(PE_101_io_data_0_out_valid),
    .io_data_0_out_bits(PE_101_io_data_0_out_bits),
    .io_sig_stat2trans(PE_101_io_sig_stat2trans)
  );
  PE PE_102 ( // @[pearray.scala 103:13]
    .clock(PE_102_clock),
    .reset(PE_102_reset),
    .io_data_2_in_valid(PE_102_io_data_2_in_valid),
    .io_data_2_in_bits(PE_102_io_data_2_in_bits),
    .io_data_2_out_valid(PE_102_io_data_2_out_valid),
    .io_data_2_out_bits(PE_102_io_data_2_out_bits),
    .io_data_1_in_valid(PE_102_io_data_1_in_valid),
    .io_data_1_in_bits(PE_102_io_data_1_in_bits),
    .io_data_1_out_valid(PE_102_io_data_1_out_valid),
    .io_data_1_out_bits(PE_102_io_data_1_out_bits),
    .io_data_0_in_valid(PE_102_io_data_0_in_valid),
    .io_data_0_in_bits(PE_102_io_data_0_in_bits),
    .io_data_0_out_valid(PE_102_io_data_0_out_valid),
    .io_data_0_out_bits(PE_102_io_data_0_out_bits),
    .io_sig_stat2trans(PE_102_io_sig_stat2trans)
  );
  PE PE_103 ( // @[pearray.scala 103:13]
    .clock(PE_103_clock),
    .reset(PE_103_reset),
    .io_data_2_in_valid(PE_103_io_data_2_in_valid),
    .io_data_2_in_bits(PE_103_io_data_2_in_bits),
    .io_data_2_out_valid(PE_103_io_data_2_out_valid),
    .io_data_2_out_bits(PE_103_io_data_2_out_bits),
    .io_data_1_in_valid(PE_103_io_data_1_in_valid),
    .io_data_1_in_bits(PE_103_io_data_1_in_bits),
    .io_data_1_out_valid(PE_103_io_data_1_out_valid),
    .io_data_1_out_bits(PE_103_io_data_1_out_bits),
    .io_data_0_in_valid(PE_103_io_data_0_in_valid),
    .io_data_0_in_bits(PE_103_io_data_0_in_bits),
    .io_data_0_out_valid(PE_103_io_data_0_out_valid),
    .io_data_0_out_bits(PE_103_io_data_0_out_bits),
    .io_sig_stat2trans(PE_103_io_sig_stat2trans)
  );
  PE PE_104 ( // @[pearray.scala 103:13]
    .clock(PE_104_clock),
    .reset(PE_104_reset),
    .io_data_2_in_valid(PE_104_io_data_2_in_valid),
    .io_data_2_in_bits(PE_104_io_data_2_in_bits),
    .io_data_2_out_valid(PE_104_io_data_2_out_valid),
    .io_data_2_out_bits(PE_104_io_data_2_out_bits),
    .io_data_1_in_valid(PE_104_io_data_1_in_valid),
    .io_data_1_in_bits(PE_104_io_data_1_in_bits),
    .io_data_1_out_valid(PE_104_io_data_1_out_valid),
    .io_data_1_out_bits(PE_104_io_data_1_out_bits),
    .io_data_0_in_valid(PE_104_io_data_0_in_valid),
    .io_data_0_in_bits(PE_104_io_data_0_in_bits),
    .io_data_0_out_valid(PE_104_io_data_0_out_valid),
    .io_data_0_out_bits(PE_104_io_data_0_out_bits),
    .io_sig_stat2trans(PE_104_io_sig_stat2trans)
  );
  PE PE_105 ( // @[pearray.scala 103:13]
    .clock(PE_105_clock),
    .reset(PE_105_reset),
    .io_data_2_in_valid(PE_105_io_data_2_in_valid),
    .io_data_2_in_bits(PE_105_io_data_2_in_bits),
    .io_data_2_out_valid(PE_105_io_data_2_out_valid),
    .io_data_2_out_bits(PE_105_io_data_2_out_bits),
    .io_data_1_in_valid(PE_105_io_data_1_in_valid),
    .io_data_1_in_bits(PE_105_io_data_1_in_bits),
    .io_data_1_out_valid(PE_105_io_data_1_out_valid),
    .io_data_1_out_bits(PE_105_io_data_1_out_bits),
    .io_data_0_in_valid(PE_105_io_data_0_in_valid),
    .io_data_0_in_bits(PE_105_io_data_0_in_bits),
    .io_data_0_out_valid(PE_105_io_data_0_out_valid),
    .io_data_0_out_bits(PE_105_io_data_0_out_bits),
    .io_sig_stat2trans(PE_105_io_sig_stat2trans)
  );
  PE PE_106 ( // @[pearray.scala 103:13]
    .clock(PE_106_clock),
    .reset(PE_106_reset),
    .io_data_2_in_valid(PE_106_io_data_2_in_valid),
    .io_data_2_in_bits(PE_106_io_data_2_in_bits),
    .io_data_2_out_valid(PE_106_io_data_2_out_valid),
    .io_data_2_out_bits(PE_106_io_data_2_out_bits),
    .io_data_1_in_valid(PE_106_io_data_1_in_valid),
    .io_data_1_in_bits(PE_106_io_data_1_in_bits),
    .io_data_1_out_valid(PE_106_io_data_1_out_valid),
    .io_data_1_out_bits(PE_106_io_data_1_out_bits),
    .io_data_0_in_valid(PE_106_io_data_0_in_valid),
    .io_data_0_in_bits(PE_106_io_data_0_in_bits),
    .io_data_0_out_valid(PE_106_io_data_0_out_valid),
    .io_data_0_out_bits(PE_106_io_data_0_out_bits),
    .io_sig_stat2trans(PE_106_io_sig_stat2trans)
  );
  PE PE_107 ( // @[pearray.scala 103:13]
    .clock(PE_107_clock),
    .reset(PE_107_reset),
    .io_data_2_in_valid(PE_107_io_data_2_in_valid),
    .io_data_2_in_bits(PE_107_io_data_2_in_bits),
    .io_data_2_out_valid(PE_107_io_data_2_out_valid),
    .io_data_2_out_bits(PE_107_io_data_2_out_bits),
    .io_data_1_in_valid(PE_107_io_data_1_in_valid),
    .io_data_1_in_bits(PE_107_io_data_1_in_bits),
    .io_data_1_out_valid(PE_107_io_data_1_out_valid),
    .io_data_1_out_bits(PE_107_io_data_1_out_bits),
    .io_data_0_in_valid(PE_107_io_data_0_in_valid),
    .io_data_0_in_bits(PE_107_io_data_0_in_bits),
    .io_data_0_out_valid(PE_107_io_data_0_out_valid),
    .io_data_0_out_bits(PE_107_io_data_0_out_bits),
    .io_sig_stat2trans(PE_107_io_sig_stat2trans)
  );
  PE PE_108 ( // @[pearray.scala 103:13]
    .clock(PE_108_clock),
    .reset(PE_108_reset),
    .io_data_2_in_valid(PE_108_io_data_2_in_valid),
    .io_data_2_in_bits(PE_108_io_data_2_in_bits),
    .io_data_2_out_valid(PE_108_io_data_2_out_valid),
    .io_data_2_out_bits(PE_108_io_data_2_out_bits),
    .io_data_1_in_valid(PE_108_io_data_1_in_valid),
    .io_data_1_in_bits(PE_108_io_data_1_in_bits),
    .io_data_1_out_valid(PE_108_io_data_1_out_valid),
    .io_data_1_out_bits(PE_108_io_data_1_out_bits),
    .io_data_0_in_valid(PE_108_io_data_0_in_valid),
    .io_data_0_in_bits(PE_108_io_data_0_in_bits),
    .io_data_0_out_valid(PE_108_io_data_0_out_valid),
    .io_data_0_out_bits(PE_108_io_data_0_out_bits),
    .io_sig_stat2trans(PE_108_io_sig_stat2trans)
  );
  PE PE_109 ( // @[pearray.scala 103:13]
    .clock(PE_109_clock),
    .reset(PE_109_reset),
    .io_data_2_in_valid(PE_109_io_data_2_in_valid),
    .io_data_2_in_bits(PE_109_io_data_2_in_bits),
    .io_data_2_out_valid(PE_109_io_data_2_out_valid),
    .io_data_2_out_bits(PE_109_io_data_2_out_bits),
    .io_data_1_in_valid(PE_109_io_data_1_in_valid),
    .io_data_1_in_bits(PE_109_io_data_1_in_bits),
    .io_data_1_out_valid(PE_109_io_data_1_out_valid),
    .io_data_1_out_bits(PE_109_io_data_1_out_bits),
    .io_data_0_in_valid(PE_109_io_data_0_in_valid),
    .io_data_0_in_bits(PE_109_io_data_0_in_bits),
    .io_data_0_out_valid(PE_109_io_data_0_out_valid),
    .io_data_0_out_bits(PE_109_io_data_0_out_bits),
    .io_sig_stat2trans(PE_109_io_sig_stat2trans)
  );
  PE PE_110 ( // @[pearray.scala 103:13]
    .clock(PE_110_clock),
    .reset(PE_110_reset),
    .io_data_2_in_valid(PE_110_io_data_2_in_valid),
    .io_data_2_in_bits(PE_110_io_data_2_in_bits),
    .io_data_2_out_valid(PE_110_io_data_2_out_valid),
    .io_data_2_out_bits(PE_110_io_data_2_out_bits),
    .io_data_1_in_valid(PE_110_io_data_1_in_valid),
    .io_data_1_in_bits(PE_110_io_data_1_in_bits),
    .io_data_1_out_valid(PE_110_io_data_1_out_valid),
    .io_data_1_out_bits(PE_110_io_data_1_out_bits),
    .io_data_0_in_valid(PE_110_io_data_0_in_valid),
    .io_data_0_in_bits(PE_110_io_data_0_in_bits),
    .io_data_0_out_valid(PE_110_io_data_0_out_valid),
    .io_data_0_out_bits(PE_110_io_data_0_out_bits),
    .io_sig_stat2trans(PE_110_io_sig_stat2trans)
  );
  PE PE_111 ( // @[pearray.scala 103:13]
    .clock(PE_111_clock),
    .reset(PE_111_reset),
    .io_data_2_in_valid(PE_111_io_data_2_in_valid),
    .io_data_2_in_bits(PE_111_io_data_2_in_bits),
    .io_data_2_out_valid(PE_111_io_data_2_out_valid),
    .io_data_2_out_bits(PE_111_io_data_2_out_bits),
    .io_data_1_in_valid(PE_111_io_data_1_in_valid),
    .io_data_1_in_bits(PE_111_io_data_1_in_bits),
    .io_data_1_out_valid(PE_111_io_data_1_out_valid),
    .io_data_1_out_bits(PE_111_io_data_1_out_bits),
    .io_data_0_in_valid(PE_111_io_data_0_in_valid),
    .io_data_0_in_bits(PE_111_io_data_0_in_bits),
    .io_data_0_out_valid(PE_111_io_data_0_out_valid),
    .io_data_0_out_bits(PE_111_io_data_0_out_bits),
    .io_sig_stat2trans(PE_111_io_sig_stat2trans)
  );
  PE PE_112 ( // @[pearray.scala 103:13]
    .clock(PE_112_clock),
    .reset(PE_112_reset),
    .io_data_2_in_valid(PE_112_io_data_2_in_valid),
    .io_data_2_in_bits(PE_112_io_data_2_in_bits),
    .io_data_2_out_valid(PE_112_io_data_2_out_valid),
    .io_data_2_out_bits(PE_112_io_data_2_out_bits),
    .io_data_1_in_valid(PE_112_io_data_1_in_valid),
    .io_data_1_in_bits(PE_112_io_data_1_in_bits),
    .io_data_1_out_valid(PE_112_io_data_1_out_valid),
    .io_data_1_out_bits(PE_112_io_data_1_out_bits),
    .io_data_0_in_valid(PE_112_io_data_0_in_valid),
    .io_data_0_in_bits(PE_112_io_data_0_in_bits),
    .io_data_0_out_valid(PE_112_io_data_0_out_valid),
    .io_data_0_out_bits(PE_112_io_data_0_out_bits),
    .io_sig_stat2trans(PE_112_io_sig_stat2trans)
  );
  PE PE_113 ( // @[pearray.scala 103:13]
    .clock(PE_113_clock),
    .reset(PE_113_reset),
    .io_data_2_in_valid(PE_113_io_data_2_in_valid),
    .io_data_2_in_bits(PE_113_io_data_2_in_bits),
    .io_data_2_out_valid(PE_113_io_data_2_out_valid),
    .io_data_2_out_bits(PE_113_io_data_2_out_bits),
    .io_data_1_in_valid(PE_113_io_data_1_in_valid),
    .io_data_1_in_bits(PE_113_io_data_1_in_bits),
    .io_data_1_out_valid(PE_113_io_data_1_out_valid),
    .io_data_1_out_bits(PE_113_io_data_1_out_bits),
    .io_data_0_in_valid(PE_113_io_data_0_in_valid),
    .io_data_0_in_bits(PE_113_io_data_0_in_bits),
    .io_data_0_out_valid(PE_113_io_data_0_out_valid),
    .io_data_0_out_bits(PE_113_io_data_0_out_bits),
    .io_sig_stat2trans(PE_113_io_sig_stat2trans)
  );
  PE PE_114 ( // @[pearray.scala 103:13]
    .clock(PE_114_clock),
    .reset(PE_114_reset),
    .io_data_2_in_valid(PE_114_io_data_2_in_valid),
    .io_data_2_in_bits(PE_114_io_data_2_in_bits),
    .io_data_2_out_valid(PE_114_io_data_2_out_valid),
    .io_data_2_out_bits(PE_114_io_data_2_out_bits),
    .io_data_1_in_valid(PE_114_io_data_1_in_valid),
    .io_data_1_in_bits(PE_114_io_data_1_in_bits),
    .io_data_1_out_valid(PE_114_io_data_1_out_valid),
    .io_data_1_out_bits(PE_114_io_data_1_out_bits),
    .io_data_0_in_valid(PE_114_io_data_0_in_valid),
    .io_data_0_in_bits(PE_114_io_data_0_in_bits),
    .io_data_0_out_valid(PE_114_io_data_0_out_valid),
    .io_data_0_out_bits(PE_114_io_data_0_out_bits),
    .io_sig_stat2trans(PE_114_io_sig_stat2trans)
  );
  PE PE_115 ( // @[pearray.scala 103:13]
    .clock(PE_115_clock),
    .reset(PE_115_reset),
    .io_data_2_in_valid(PE_115_io_data_2_in_valid),
    .io_data_2_in_bits(PE_115_io_data_2_in_bits),
    .io_data_2_out_valid(PE_115_io_data_2_out_valid),
    .io_data_2_out_bits(PE_115_io_data_2_out_bits),
    .io_data_1_in_valid(PE_115_io_data_1_in_valid),
    .io_data_1_in_bits(PE_115_io_data_1_in_bits),
    .io_data_1_out_valid(PE_115_io_data_1_out_valid),
    .io_data_1_out_bits(PE_115_io_data_1_out_bits),
    .io_data_0_in_valid(PE_115_io_data_0_in_valid),
    .io_data_0_in_bits(PE_115_io_data_0_in_bits),
    .io_data_0_out_valid(PE_115_io_data_0_out_valid),
    .io_data_0_out_bits(PE_115_io_data_0_out_bits),
    .io_sig_stat2trans(PE_115_io_sig_stat2trans)
  );
  PE PE_116 ( // @[pearray.scala 103:13]
    .clock(PE_116_clock),
    .reset(PE_116_reset),
    .io_data_2_in_valid(PE_116_io_data_2_in_valid),
    .io_data_2_in_bits(PE_116_io_data_2_in_bits),
    .io_data_2_out_valid(PE_116_io_data_2_out_valid),
    .io_data_2_out_bits(PE_116_io_data_2_out_bits),
    .io_data_1_in_valid(PE_116_io_data_1_in_valid),
    .io_data_1_in_bits(PE_116_io_data_1_in_bits),
    .io_data_1_out_valid(PE_116_io_data_1_out_valid),
    .io_data_1_out_bits(PE_116_io_data_1_out_bits),
    .io_data_0_in_valid(PE_116_io_data_0_in_valid),
    .io_data_0_in_bits(PE_116_io_data_0_in_bits),
    .io_data_0_out_valid(PE_116_io_data_0_out_valid),
    .io_data_0_out_bits(PE_116_io_data_0_out_bits),
    .io_sig_stat2trans(PE_116_io_sig_stat2trans)
  );
  PE PE_117 ( // @[pearray.scala 103:13]
    .clock(PE_117_clock),
    .reset(PE_117_reset),
    .io_data_2_in_valid(PE_117_io_data_2_in_valid),
    .io_data_2_in_bits(PE_117_io_data_2_in_bits),
    .io_data_2_out_valid(PE_117_io_data_2_out_valid),
    .io_data_2_out_bits(PE_117_io_data_2_out_bits),
    .io_data_1_in_valid(PE_117_io_data_1_in_valid),
    .io_data_1_in_bits(PE_117_io_data_1_in_bits),
    .io_data_1_out_valid(PE_117_io_data_1_out_valid),
    .io_data_1_out_bits(PE_117_io_data_1_out_bits),
    .io_data_0_in_valid(PE_117_io_data_0_in_valid),
    .io_data_0_in_bits(PE_117_io_data_0_in_bits),
    .io_data_0_out_valid(PE_117_io_data_0_out_valid),
    .io_data_0_out_bits(PE_117_io_data_0_out_bits),
    .io_sig_stat2trans(PE_117_io_sig_stat2trans)
  );
  PE PE_118 ( // @[pearray.scala 103:13]
    .clock(PE_118_clock),
    .reset(PE_118_reset),
    .io_data_2_in_valid(PE_118_io_data_2_in_valid),
    .io_data_2_in_bits(PE_118_io_data_2_in_bits),
    .io_data_2_out_valid(PE_118_io_data_2_out_valid),
    .io_data_2_out_bits(PE_118_io_data_2_out_bits),
    .io_data_1_in_valid(PE_118_io_data_1_in_valid),
    .io_data_1_in_bits(PE_118_io_data_1_in_bits),
    .io_data_1_out_valid(PE_118_io_data_1_out_valid),
    .io_data_1_out_bits(PE_118_io_data_1_out_bits),
    .io_data_0_in_valid(PE_118_io_data_0_in_valid),
    .io_data_0_in_bits(PE_118_io_data_0_in_bits),
    .io_data_0_out_valid(PE_118_io_data_0_out_valid),
    .io_data_0_out_bits(PE_118_io_data_0_out_bits),
    .io_sig_stat2trans(PE_118_io_sig_stat2trans)
  );
  PE PE_119 ( // @[pearray.scala 103:13]
    .clock(PE_119_clock),
    .reset(PE_119_reset),
    .io_data_2_in_valid(PE_119_io_data_2_in_valid),
    .io_data_2_in_bits(PE_119_io_data_2_in_bits),
    .io_data_2_out_valid(PE_119_io_data_2_out_valid),
    .io_data_2_out_bits(PE_119_io_data_2_out_bits),
    .io_data_1_in_valid(PE_119_io_data_1_in_valid),
    .io_data_1_in_bits(PE_119_io_data_1_in_bits),
    .io_data_1_out_valid(PE_119_io_data_1_out_valid),
    .io_data_1_out_bits(PE_119_io_data_1_out_bits),
    .io_data_0_in_valid(PE_119_io_data_0_in_valid),
    .io_data_0_in_bits(PE_119_io_data_0_in_bits),
    .io_data_0_out_valid(PE_119_io_data_0_out_valid),
    .io_data_0_out_bits(PE_119_io_data_0_out_bits),
    .io_sig_stat2trans(PE_119_io_sig_stat2trans)
  );
  PE PE_120 ( // @[pearray.scala 103:13]
    .clock(PE_120_clock),
    .reset(PE_120_reset),
    .io_data_2_in_valid(PE_120_io_data_2_in_valid),
    .io_data_2_in_bits(PE_120_io_data_2_in_bits),
    .io_data_2_out_valid(PE_120_io_data_2_out_valid),
    .io_data_2_out_bits(PE_120_io_data_2_out_bits),
    .io_data_1_in_valid(PE_120_io_data_1_in_valid),
    .io_data_1_in_bits(PE_120_io_data_1_in_bits),
    .io_data_1_out_valid(PE_120_io_data_1_out_valid),
    .io_data_1_out_bits(PE_120_io_data_1_out_bits),
    .io_data_0_in_valid(PE_120_io_data_0_in_valid),
    .io_data_0_in_bits(PE_120_io_data_0_in_bits),
    .io_data_0_out_valid(PE_120_io_data_0_out_valid),
    .io_data_0_out_bits(PE_120_io_data_0_out_bits),
    .io_sig_stat2trans(PE_120_io_sig_stat2trans)
  );
  PE PE_121 ( // @[pearray.scala 103:13]
    .clock(PE_121_clock),
    .reset(PE_121_reset),
    .io_data_2_in_valid(PE_121_io_data_2_in_valid),
    .io_data_2_in_bits(PE_121_io_data_2_in_bits),
    .io_data_2_out_valid(PE_121_io_data_2_out_valid),
    .io_data_2_out_bits(PE_121_io_data_2_out_bits),
    .io_data_1_in_valid(PE_121_io_data_1_in_valid),
    .io_data_1_in_bits(PE_121_io_data_1_in_bits),
    .io_data_1_out_valid(PE_121_io_data_1_out_valid),
    .io_data_1_out_bits(PE_121_io_data_1_out_bits),
    .io_data_0_in_valid(PE_121_io_data_0_in_valid),
    .io_data_0_in_bits(PE_121_io_data_0_in_bits),
    .io_data_0_out_valid(PE_121_io_data_0_out_valid),
    .io_data_0_out_bits(PE_121_io_data_0_out_bits),
    .io_sig_stat2trans(PE_121_io_sig_stat2trans)
  );
  PE PE_122 ( // @[pearray.scala 103:13]
    .clock(PE_122_clock),
    .reset(PE_122_reset),
    .io_data_2_in_valid(PE_122_io_data_2_in_valid),
    .io_data_2_in_bits(PE_122_io_data_2_in_bits),
    .io_data_2_out_valid(PE_122_io_data_2_out_valid),
    .io_data_2_out_bits(PE_122_io_data_2_out_bits),
    .io_data_1_in_valid(PE_122_io_data_1_in_valid),
    .io_data_1_in_bits(PE_122_io_data_1_in_bits),
    .io_data_1_out_valid(PE_122_io_data_1_out_valid),
    .io_data_1_out_bits(PE_122_io_data_1_out_bits),
    .io_data_0_in_valid(PE_122_io_data_0_in_valid),
    .io_data_0_in_bits(PE_122_io_data_0_in_bits),
    .io_data_0_out_valid(PE_122_io_data_0_out_valid),
    .io_data_0_out_bits(PE_122_io_data_0_out_bits),
    .io_sig_stat2trans(PE_122_io_sig_stat2trans)
  );
  PE PE_123 ( // @[pearray.scala 103:13]
    .clock(PE_123_clock),
    .reset(PE_123_reset),
    .io_data_2_in_valid(PE_123_io_data_2_in_valid),
    .io_data_2_in_bits(PE_123_io_data_2_in_bits),
    .io_data_2_out_valid(PE_123_io_data_2_out_valid),
    .io_data_2_out_bits(PE_123_io_data_2_out_bits),
    .io_data_1_in_valid(PE_123_io_data_1_in_valid),
    .io_data_1_in_bits(PE_123_io_data_1_in_bits),
    .io_data_1_out_valid(PE_123_io_data_1_out_valid),
    .io_data_1_out_bits(PE_123_io_data_1_out_bits),
    .io_data_0_in_valid(PE_123_io_data_0_in_valid),
    .io_data_0_in_bits(PE_123_io_data_0_in_bits),
    .io_data_0_out_valid(PE_123_io_data_0_out_valid),
    .io_data_0_out_bits(PE_123_io_data_0_out_bits),
    .io_sig_stat2trans(PE_123_io_sig_stat2trans)
  );
  PE PE_124 ( // @[pearray.scala 103:13]
    .clock(PE_124_clock),
    .reset(PE_124_reset),
    .io_data_2_in_valid(PE_124_io_data_2_in_valid),
    .io_data_2_in_bits(PE_124_io_data_2_in_bits),
    .io_data_2_out_valid(PE_124_io_data_2_out_valid),
    .io_data_2_out_bits(PE_124_io_data_2_out_bits),
    .io_data_1_in_valid(PE_124_io_data_1_in_valid),
    .io_data_1_in_bits(PE_124_io_data_1_in_bits),
    .io_data_1_out_valid(PE_124_io_data_1_out_valid),
    .io_data_1_out_bits(PE_124_io_data_1_out_bits),
    .io_data_0_in_valid(PE_124_io_data_0_in_valid),
    .io_data_0_in_bits(PE_124_io_data_0_in_bits),
    .io_data_0_out_valid(PE_124_io_data_0_out_valid),
    .io_data_0_out_bits(PE_124_io_data_0_out_bits),
    .io_sig_stat2trans(PE_124_io_sig_stat2trans)
  );
  PE PE_125 ( // @[pearray.scala 103:13]
    .clock(PE_125_clock),
    .reset(PE_125_reset),
    .io_data_2_in_valid(PE_125_io_data_2_in_valid),
    .io_data_2_in_bits(PE_125_io_data_2_in_bits),
    .io_data_2_out_valid(PE_125_io_data_2_out_valid),
    .io_data_2_out_bits(PE_125_io_data_2_out_bits),
    .io_data_1_in_valid(PE_125_io_data_1_in_valid),
    .io_data_1_in_bits(PE_125_io_data_1_in_bits),
    .io_data_1_out_valid(PE_125_io_data_1_out_valid),
    .io_data_1_out_bits(PE_125_io_data_1_out_bits),
    .io_data_0_in_valid(PE_125_io_data_0_in_valid),
    .io_data_0_in_bits(PE_125_io_data_0_in_bits),
    .io_data_0_out_valid(PE_125_io_data_0_out_valid),
    .io_data_0_out_bits(PE_125_io_data_0_out_bits),
    .io_sig_stat2trans(PE_125_io_sig_stat2trans)
  );
  PE PE_126 ( // @[pearray.scala 103:13]
    .clock(PE_126_clock),
    .reset(PE_126_reset),
    .io_data_2_in_valid(PE_126_io_data_2_in_valid),
    .io_data_2_in_bits(PE_126_io_data_2_in_bits),
    .io_data_2_out_valid(PE_126_io_data_2_out_valid),
    .io_data_2_out_bits(PE_126_io_data_2_out_bits),
    .io_data_1_in_valid(PE_126_io_data_1_in_valid),
    .io_data_1_in_bits(PE_126_io_data_1_in_bits),
    .io_data_1_out_valid(PE_126_io_data_1_out_valid),
    .io_data_1_out_bits(PE_126_io_data_1_out_bits),
    .io_data_0_in_valid(PE_126_io_data_0_in_valid),
    .io_data_0_in_bits(PE_126_io_data_0_in_bits),
    .io_data_0_out_valid(PE_126_io_data_0_out_valid),
    .io_data_0_out_bits(PE_126_io_data_0_out_bits),
    .io_sig_stat2trans(PE_126_io_sig_stat2trans)
  );
  PE PE_127 ( // @[pearray.scala 103:13]
    .clock(PE_127_clock),
    .reset(PE_127_reset),
    .io_data_2_in_valid(PE_127_io_data_2_in_valid),
    .io_data_2_in_bits(PE_127_io_data_2_in_bits),
    .io_data_2_out_valid(PE_127_io_data_2_out_valid),
    .io_data_2_out_bits(PE_127_io_data_2_out_bits),
    .io_data_1_in_valid(PE_127_io_data_1_in_valid),
    .io_data_1_in_bits(PE_127_io_data_1_in_bits),
    .io_data_1_out_valid(PE_127_io_data_1_out_valid),
    .io_data_1_out_bits(PE_127_io_data_1_out_bits),
    .io_data_0_in_valid(PE_127_io_data_0_in_valid),
    .io_data_0_in_bits(PE_127_io_data_0_in_bits),
    .io_data_0_out_valid(PE_127_io_data_0_out_valid),
    .io_data_0_out_bits(PE_127_io_data_0_out_bits),
    .io_sig_stat2trans(PE_127_io_sig_stat2trans)
  );
  PE PE_128 ( // @[pearray.scala 103:13]
    .clock(PE_128_clock),
    .reset(PE_128_reset),
    .io_data_2_in_valid(PE_128_io_data_2_in_valid),
    .io_data_2_in_bits(PE_128_io_data_2_in_bits),
    .io_data_2_out_valid(PE_128_io_data_2_out_valid),
    .io_data_2_out_bits(PE_128_io_data_2_out_bits),
    .io_data_1_in_valid(PE_128_io_data_1_in_valid),
    .io_data_1_in_bits(PE_128_io_data_1_in_bits),
    .io_data_1_out_valid(PE_128_io_data_1_out_valid),
    .io_data_1_out_bits(PE_128_io_data_1_out_bits),
    .io_data_0_in_valid(PE_128_io_data_0_in_valid),
    .io_data_0_in_bits(PE_128_io_data_0_in_bits),
    .io_data_0_out_valid(PE_128_io_data_0_out_valid),
    .io_data_0_out_bits(PE_128_io_data_0_out_bits),
    .io_sig_stat2trans(PE_128_io_sig_stat2trans)
  );
  PE PE_129 ( // @[pearray.scala 103:13]
    .clock(PE_129_clock),
    .reset(PE_129_reset),
    .io_data_2_in_valid(PE_129_io_data_2_in_valid),
    .io_data_2_in_bits(PE_129_io_data_2_in_bits),
    .io_data_2_out_valid(PE_129_io_data_2_out_valid),
    .io_data_2_out_bits(PE_129_io_data_2_out_bits),
    .io_data_1_in_valid(PE_129_io_data_1_in_valid),
    .io_data_1_in_bits(PE_129_io_data_1_in_bits),
    .io_data_1_out_valid(PE_129_io_data_1_out_valid),
    .io_data_1_out_bits(PE_129_io_data_1_out_bits),
    .io_data_0_in_valid(PE_129_io_data_0_in_valid),
    .io_data_0_in_bits(PE_129_io_data_0_in_bits),
    .io_data_0_out_valid(PE_129_io_data_0_out_valid),
    .io_data_0_out_bits(PE_129_io_data_0_out_bits),
    .io_sig_stat2trans(PE_129_io_sig_stat2trans)
  );
  PE PE_130 ( // @[pearray.scala 103:13]
    .clock(PE_130_clock),
    .reset(PE_130_reset),
    .io_data_2_in_valid(PE_130_io_data_2_in_valid),
    .io_data_2_in_bits(PE_130_io_data_2_in_bits),
    .io_data_2_out_valid(PE_130_io_data_2_out_valid),
    .io_data_2_out_bits(PE_130_io_data_2_out_bits),
    .io_data_1_in_valid(PE_130_io_data_1_in_valid),
    .io_data_1_in_bits(PE_130_io_data_1_in_bits),
    .io_data_1_out_valid(PE_130_io_data_1_out_valid),
    .io_data_1_out_bits(PE_130_io_data_1_out_bits),
    .io_data_0_in_valid(PE_130_io_data_0_in_valid),
    .io_data_0_in_bits(PE_130_io_data_0_in_bits),
    .io_data_0_out_valid(PE_130_io_data_0_out_valid),
    .io_data_0_out_bits(PE_130_io_data_0_out_bits),
    .io_sig_stat2trans(PE_130_io_sig_stat2trans)
  );
  PE PE_131 ( // @[pearray.scala 103:13]
    .clock(PE_131_clock),
    .reset(PE_131_reset),
    .io_data_2_in_valid(PE_131_io_data_2_in_valid),
    .io_data_2_in_bits(PE_131_io_data_2_in_bits),
    .io_data_2_out_valid(PE_131_io_data_2_out_valid),
    .io_data_2_out_bits(PE_131_io_data_2_out_bits),
    .io_data_1_in_valid(PE_131_io_data_1_in_valid),
    .io_data_1_in_bits(PE_131_io_data_1_in_bits),
    .io_data_1_out_valid(PE_131_io_data_1_out_valid),
    .io_data_1_out_bits(PE_131_io_data_1_out_bits),
    .io_data_0_in_valid(PE_131_io_data_0_in_valid),
    .io_data_0_in_bits(PE_131_io_data_0_in_bits),
    .io_data_0_out_valid(PE_131_io_data_0_out_valid),
    .io_data_0_out_bits(PE_131_io_data_0_out_bits),
    .io_sig_stat2trans(PE_131_io_sig_stat2trans)
  );
  PE PE_132 ( // @[pearray.scala 103:13]
    .clock(PE_132_clock),
    .reset(PE_132_reset),
    .io_data_2_in_valid(PE_132_io_data_2_in_valid),
    .io_data_2_in_bits(PE_132_io_data_2_in_bits),
    .io_data_2_out_valid(PE_132_io_data_2_out_valid),
    .io_data_2_out_bits(PE_132_io_data_2_out_bits),
    .io_data_1_in_valid(PE_132_io_data_1_in_valid),
    .io_data_1_in_bits(PE_132_io_data_1_in_bits),
    .io_data_1_out_valid(PE_132_io_data_1_out_valid),
    .io_data_1_out_bits(PE_132_io_data_1_out_bits),
    .io_data_0_in_valid(PE_132_io_data_0_in_valid),
    .io_data_0_in_bits(PE_132_io_data_0_in_bits),
    .io_data_0_out_valid(PE_132_io_data_0_out_valid),
    .io_data_0_out_bits(PE_132_io_data_0_out_bits),
    .io_sig_stat2trans(PE_132_io_sig_stat2trans)
  );
  PE PE_133 ( // @[pearray.scala 103:13]
    .clock(PE_133_clock),
    .reset(PE_133_reset),
    .io_data_2_in_valid(PE_133_io_data_2_in_valid),
    .io_data_2_in_bits(PE_133_io_data_2_in_bits),
    .io_data_2_out_valid(PE_133_io_data_2_out_valid),
    .io_data_2_out_bits(PE_133_io_data_2_out_bits),
    .io_data_1_in_valid(PE_133_io_data_1_in_valid),
    .io_data_1_in_bits(PE_133_io_data_1_in_bits),
    .io_data_1_out_valid(PE_133_io_data_1_out_valid),
    .io_data_1_out_bits(PE_133_io_data_1_out_bits),
    .io_data_0_in_valid(PE_133_io_data_0_in_valid),
    .io_data_0_in_bits(PE_133_io_data_0_in_bits),
    .io_data_0_out_valid(PE_133_io_data_0_out_valid),
    .io_data_0_out_bits(PE_133_io_data_0_out_bits),
    .io_sig_stat2trans(PE_133_io_sig_stat2trans)
  );
  PE PE_134 ( // @[pearray.scala 103:13]
    .clock(PE_134_clock),
    .reset(PE_134_reset),
    .io_data_2_in_valid(PE_134_io_data_2_in_valid),
    .io_data_2_in_bits(PE_134_io_data_2_in_bits),
    .io_data_2_out_valid(PE_134_io_data_2_out_valid),
    .io_data_2_out_bits(PE_134_io_data_2_out_bits),
    .io_data_1_in_valid(PE_134_io_data_1_in_valid),
    .io_data_1_in_bits(PE_134_io_data_1_in_bits),
    .io_data_1_out_valid(PE_134_io_data_1_out_valid),
    .io_data_1_out_bits(PE_134_io_data_1_out_bits),
    .io_data_0_in_valid(PE_134_io_data_0_in_valid),
    .io_data_0_in_bits(PE_134_io_data_0_in_bits),
    .io_data_0_out_valid(PE_134_io_data_0_out_valid),
    .io_data_0_out_bits(PE_134_io_data_0_out_bits),
    .io_sig_stat2trans(PE_134_io_sig_stat2trans)
  );
  PE PE_135 ( // @[pearray.scala 103:13]
    .clock(PE_135_clock),
    .reset(PE_135_reset),
    .io_data_2_in_valid(PE_135_io_data_2_in_valid),
    .io_data_2_in_bits(PE_135_io_data_2_in_bits),
    .io_data_2_out_valid(PE_135_io_data_2_out_valid),
    .io_data_2_out_bits(PE_135_io_data_2_out_bits),
    .io_data_1_in_valid(PE_135_io_data_1_in_valid),
    .io_data_1_in_bits(PE_135_io_data_1_in_bits),
    .io_data_1_out_valid(PE_135_io_data_1_out_valid),
    .io_data_1_out_bits(PE_135_io_data_1_out_bits),
    .io_data_0_in_valid(PE_135_io_data_0_in_valid),
    .io_data_0_in_bits(PE_135_io_data_0_in_bits),
    .io_data_0_out_valid(PE_135_io_data_0_out_valid),
    .io_data_0_out_bits(PE_135_io_data_0_out_bits),
    .io_sig_stat2trans(PE_135_io_sig_stat2trans)
  );
  PE PE_136 ( // @[pearray.scala 103:13]
    .clock(PE_136_clock),
    .reset(PE_136_reset),
    .io_data_2_in_valid(PE_136_io_data_2_in_valid),
    .io_data_2_in_bits(PE_136_io_data_2_in_bits),
    .io_data_2_out_valid(PE_136_io_data_2_out_valid),
    .io_data_2_out_bits(PE_136_io_data_2_out_bits),
    .io_data_1_in_valid(PE_136_io_data_1_in_valid),
    .io_data_1_in_bits(PE_136_io_data_1_in_bits),
    .io_data_1_out_valid(PE_136_io_data_1_out_valid),
    .io_data_1_out_bits(PE_136_io_data_1_out_bits),
    .io_data_0_in_valid(PE_136_io_data_0_in_valid),
    .io_data_0_in_bits(PE_136_io_data_0_in_bits),
    .io_data_0_out_valid(PE_136_io_data_0_out_valid),
    .io_data_0_out_bits(PE_136_io_data_0_out_bits),
    .io_sig_stat2trans(PE_136_io_sig_stat2trans)
  );
  PE PE_137 ( // @[pearray.scala 103:13]
    .clock(PE_137_clock),
    .reset(PE_137_reset),
    .io_data_2_in_valid(PE_137_io_data_2_in_valid),
    .io_data_2_in_bits(PE_137_io_data_2_in_bits),
    .io_data_2_out_valid(PE_137_io_data_2_out_valid),
    .io_data_2_out_bits(PE_137_io_data_2_out_bits),
    .io_data_1_in_valid(PE_137_io_data_1_in_valid),
    .io_data_1_in_bits(PE_137_io_data_1_in_bits),
    .io_data_1_out_valid(PE_137_io_data_1_out_valid),
    .io_data_1_out_bits(PE_137_io_data_1_out_bits),
    .io_data_0_in_valid(PE_137_io_data_0_in_valid),
    .io_data_0_in_bits(PE_137_io_data_0_in_bits),
    .io_data_0_out_valid(PE_137_io_data_0_out_valid),
    .io_data_0_out_bits(PE_137_io_data_0_out_bits),
    .io_sig_stat2trans(PE_137_io_sig_stat2trans)
  );
  PE PE_138 ( // @[pearray.scala 103:13]
    .clock(PE_138_clock),
    .reset(PE_138_reset),
    .io_data_2_in_valid(PE_138_io_data_2_in_valid),
    .io_data_2_in_bits(PE_138_io_data_2_in_bits),
    .io_data_2_out_valid(PE_138_io_data_2_out_valid),
    .io_data_2_out_bits(PE_138_io_data_2_out_bits),
    .io_data_1_in_valid(PE_138_io_data_1_in_valid),
    .io_data_1_in_bits(PE_138_io_data_1_in_bits),
    .io_data_1_out_valid(PE_138_io_data_1_out_valid),
    .io_data_1_out_bits(PE_138_io_data_1_out_bits),
    .io_data_0_in_valid(PE_138_io_data_0_in_valid),
    .io_data_0_in_bits(PE_138_io_data_0_in_bits),
    .io_data_0_out_valid(PE_138_io_data_0_out_valid),
    .io_data_0_out_bits(PE_138_io_data_0_out_bits),
    .io_sig_stat2trans(PE_138_io_sig_stat2trans)
  );
  PE PE_139 ( // @[pearray.scala 103:13]
    .clock(PE_139_clock),
    .reset(PE_139_reset),
    .io_data_2_in_valid(PE_139_io_data_2_in_valid),
    .io_data_2_in_bits(PE_139_io_data_2_in_bits),
    .io_data_2_out_valid(PE_139_io_data_2_out_valid),
    .io_data_2_out_bits(PE_139_io_data_2_out_bits),
    .io_data_1_in_valid(PE_139_io_data_1_in_valid),
    .io_data_1_in_bits(PE_139_io_data_1_in_bits),
    .io_data_1_out_valid(PE_139_io_data_1_out_valid),
    .io_data_1_out_bits(PE_139_io_data_1_out_bits),
    .io_data_0_in_valid(PE_139_io_data_0_in_valid),
    .io_data_0_in_bits(PE_139_io_data_0_in_bits),
    .io_data_0_out_valid(PE_139_io_data_0_out_valid),
    .io_data_0_out_bits(PE_139_io_data_0_out_bits),
    .io_sig_stat2trans(PE_139_io_sig_stat2trans)
  );
  PE PE_140 ( // @[pearray.scala 103:13]
    .clock(PE_140_clock),
    .reset(PE_140_reset),
    .io_data_2_in_valid(PE_140_io_data_2_in_valid),
    .io_data_2_in_bits(PE_140_io_data_2_in_bits),
    .io_data_2_out_valid(PE_140_io_data_2_out_valid),
    .io_data_2_out_bits(PE_140_io_data_2_out_bits),
    .io_data_1_in_valid(PE_140_io_data_1_in_valid),
    .io_data_1_in_bits(PE_140_io_data_1_in_bits),
    .io_data_1_out_valid(PE_140_io_data_1_out_valid),
    .io_data_1_out_bits(PE_140_io_data_1_out_bits),
    .io_data_0_in_valid(PE_140_io_data_0_in_valid),
    .io_data_0_in_bits(PE_140_io_data_0_in_bits),
    .io_data_0_out_valid(PE_140_io_data_0_out_valid),
    .io_data_0_out_bits(PE_140_io_data_0_out_bits),
    .io_sig_stat2trans(PE_140_io_sig_stat2trans)
  );
  PE PE_141 ( // @[pearray.scala 103:13]
    .clock(PE_141_clock),
    .reset(PE_141_reset),
    .io_data_2_in_valid(PE_141_io_data_2_in_valid),
    .io_data_2_in_bits(PE_141_io_data_2_in_bits),
    .io_data_2_out_valid(PE_141_io_data_2_out_valid),
    .io_data_2_out_bits(PE_141_io_data_2_out_bits),
    .io_data_1_in_valid(PE_141_io_data_1_in_valid),
    .io_data_1_in_bits(PE_141_io_data_1_in_bits),
    .io_data_1_out_valid(PE_141_io_data_1_out_valid),
    .io_data_1_out_bits(PE_141_io_data_1_out_bits),
    .io_data_0_in_valid(PE_141_io_data_0_in_valid),
    .io_data_0_in_bits(PE_141_io_data_0_in_bits),
    .io_data_0_out_valid(PE_141_io_data_0_out_valid),
    .io_data_0_out_bits(PE_141_io_data_0_out_bits),
    .io_sig_stat2trans(PE_141_io_sig_stat2trans)
  );
  PE PE_142 ( // @[pearray.scala 103:13]
    .clock(PE_142_clock),
    .reset(PE_142_reset),
    .io_data_2_in_valid(PE_142_io_data_2_in_valid),
    .io_data_2_in_bits(PE_142_io_data_2_in_bits),
    .io_data_2_out_valid(PE_142_io_data_2_out_valid),
    .io_data_2_out_bits(PE_142_io_data_2_out_bits),
    .io_data_1_in_valid(PE_142_io_data_1_in_valid),
    .io_data_1_in_bits(PE_142_io_data_1_in_bits),
    .io_data_1_out_valid(PE_142_io_data_1_out_valid),
    .io_data_1_out_bits(PE_142_io_data_1_out_bits),
    .io_data_0_in_valid(PE_142_io_data_0_in_valid),
    .io_data_0_in_bits(PE_142_io_data_0_in_bits),
    .io_data_0_out_valid(PE_142_io_data_0_out_valid),
    .io_data_0_out_bits(PE_142_io_data_0_out_bits),
    .io_sig_stat2trans(PE_142_io_sig_stat2trans)
  );
  PE PE_143 ( // @[pearray.scala 103:13]
    .clock(PE_143_clock),
    .reset(PE_143_reset),
    .io_data_2_in_valid(PE_143_io_data_2_in_valid),
    .io_data_2_in_bits(PE_143_io_data_2_in_bits),
    .io_data_2_out_valid(PE_143_io_data_2_out_valid),
    .io_data_2_out_bits(PE_143_io_data_2_out_bits),
    .io_data_1_in_valid(PE_143_io_data_1_in_valid),
    .io_data_1_in_bits(PE_143_io_data_1_in_bits),
    .io_data_1_out_valid(PE_143_io_data_1_out_valid),
    .io_data_1_out_bits(PE_143_io_data_1_out_bits),
    .io_data_0_in_valid(PE_143_io_data_0_in_valid),
    .io_data_0_in_bits(PE_143_io_data_0_in_bits),
    .io_data_0_out_valid(PE_143_io_data_0_out_valid),
    .io_data_0_out_bits(PE_143_io_data_0_out_bits),
    .io_sig_stat2trans(PE_143_io_sig_stat2trans)
  );
  PE PE_144 ( // @[pearray.scala 103:13]
    .clock(PE_144_clock),
    .reset(PE_144_reset),
    .io_data_2_in_valid(PE_144_io_data_2_in_valid),
    .io_data_2_in_bits(PE_144_io_data_2_in_bits),
    .io_data_2_out_valid(PE_144_io_data_2_out_valid),
    .io_data_2_out_bits(PE_144_io_data_2_out_bits),
    .io_data_1_in_valid(PE_144_io_data_1_in_valid),
    .io_data_1_in_bits(PE_144_io_data_1_in_bits),
    .io_data_1_out_valid(PE_144_io_data_1_out_valid),
    .io_data_1_out_bits(PE_144_io_data_1_out_bits),
    .io_data_0_in_valid(PE_144_io_data_0_in_valid),
    .io_data_0_in_bits(PE_144_io_data_0_in_bits),
    .io_data_0_out_valid(PE_144_io_data_0_out_valid),
    .io_data_0_out_bits(PE_144_io_data_0_out_bits),
    .io_sig_stat2trans(PE_144_io_sig_stat2trans)
  );
  PE PE_145 ( // @[pearray.scala 103:13]
    .clock(PE_145_clock),
    .reset(PE_145_reset),
    .io_data_2_in_valid(PE_145_io_data_2_in_valid),
    .io_data_2_in_bits(PE_145_io_data_2_in_bits),
    .io_data_2_out_valid(PE_145_io_data_2_out_valid),
    .io_data_2_out_bits(PE_145_io_data_2_out_bits),
    .io_data_1_in_valid(PE_145_io_data_1_in_valid),
    .io_data_1_in_bits(PE_145_io_data_1_in_bits),
    .io_data_1_out_valid(PE_145_io_data_1_out_valid),
    .io_data_1_out_bits(PE_145_io_data_1_out_bits),
    .io_data_0_in_valid(PE_145_io_data_0_in_valid),
    .io_data_0_in_bits(PE_145_io_data_0_in_bits),
    .io_data_0_out_valid(PE_145_io_data_0_out_valid),
    .io_data_0_out_bits(PE_145_io_data_0_out_bits),
    .io_sig_stat2trans(PE_145_io_sig_stat2trans)
  );
  PE PE_146 ( // @[pearray.scala 103:13]
    .clock(PE_146_clock),
    .reset(PE_146_reset),
    .io_data_2_in_valid(PE_146_io_data_2_in_valid),
    .io_data_2_in_bits(PE_146_io_data_2_in_bits),
    .io_data_2_out_valid(PE_146_io_data_2_out_valid),
    .io_data_2_out_bits(PE_146_io_data_2_out_bits),
    .io_data_1_in_valid(PE_146_io_data_1_in_valid),
    .io_data_1_in_bits(PE_146_io_data_1_in_bits),
    .io_data_1_out_valid(PE_146_io_data_1_out_valid),
    .io_data_1_out_bits(PE_146_io_data_1_out_bits),
    .io_data_0_in_valid(PE_146_io_data_0_in_valid),
    .io_data_0_in_bits(PE_146_io_data_0_in_bits),
    .io_data_0_out_valid(PE_146_io_data_0_out_valid),
    .io_data_0_out_bits(PE_146_io_data_0_out_bits),
    .io_sig_stat2trans(PE_146_io_sig_stat2trans)
  );
  PE PE_147 ( // @[pearray.scala 103:13]
    .clock(PE_147_clock),
    .reset(PE_147_reset),
    .io_data_2_in_valid(PE_147_io_data_2_in_valid),
    .io_data_2_in_bits(PE_147_io_data_2_in_bits),
    .io_data_2_out_valid(PE_147_io_data_2_out_valid),
    .io_data_2_out_bits(PE_147_io_data_2_out_bits),
    .io_data_1_in_valid(PE_147_io_data_1_in_valid),
    .io_data_1_in_bits(PE_147_io_data_1_in_bits),
    .io_data_1_out_valid(PE_147_io_data_1_out_valid),
    .io_data_1_out_bits(PE_147_io_data_1_out_bits),
    .io_data_0_in_valid(PE_147_io_data_0_in_valid),
    .io_data_0_in_bits(PE_147_io_data_0_in_bits),
    .io_data_0_out_valid(PE_147_io_data_0_out_valid),
    .io_data_0_out_bits(PE_147_io_data_0_out_bits),
    .io_sig_stat2trans(PE_147_io_sig_stat2trans)
  );
  PE PE_148 ( // @[pearray.scala 103:13]
    .clock(PE_148_clock),
    .reset(PE_148_reset),
    .io_data_2_in_valid(PE_148_io_data_2_in_valid),
    .io_data_2_in_bits(PE_148_io_data_2_in_bits),
    .io_data_2_out_valid(PE_148_io_data_2_out_valid),
    .io_data_2_out_bits(PE_148_io_data_2_out_bits),
    .io_data_1_in_valid(PE_148_io_data_1_in_valid),
    .io_data_1_in_bits(PE_148_io_data_1_in_bits),
    .io_data_1_out_valid(PE_148_io_data_1_out_valid),
    .io_data_1_out_bits(PE_148_io_data_1_out_bits),
    .io_data_0_in_valid(PE_148_io_data_0_in_valid),
    .io_data_0_in_bits(PE_148_io_data_0_in_bits),
    .io_data_0_out_valid(PE_148_io_data_0_out_valid),
    .io_data_0_out_bits(PE_148_io_data_0_out_bits),
    .io_sig_stat2trans(PE_148_io_sig_stat2trans)
  );
  PE PE_149 ( // @[pearray.scala 103:13]
    .clock(PE_149_clock),
    .reset(PE_149_reset),
    .io_data_2_in_valid(PE_149_io_data_2_in_valid),
    .io_data_2_in_bits(PE_149_io_data_2_in_bits),
    .io_data_2_out_valid(PE_149_io_data_2_out_valid),
    .io_data_2_out_bits(PE_149_io_data_2_out_bits),
    .io_data_1_in_valid(PE_149_io_data_1_in_valid),
    .io_data_1_in_bits(PE_149_io_data_1_in_bits),
    .io_data_1_out_valid(PE_149_io_data_1_out_valid),
    .io_data_1_out_bits(PE_149_io_data_1_out_bits),
    .io_data_0_in_valid(PE_149_io_data_0_in_valid),
    .io_data_0_in_bits(PE_149_io_data_0_in_bits),
    .io_data_0_out_valid(PE_149_io_data_0_out_valid),
    .io_data_0_out_bits(PE_149_io_data_0_out_bits),
    .io_sig_stat2trans(PE_149_io_sig_stat2trans)
  );
  PE PE_150 ( // @[pearray.scala 103:13]
    .clock(PE_150_clock),
    .reset(PE_150_reset),
    .io_data_2_in_valid(PE_150_io_data_2_in_valid),
    .io_data_2_in_bits(PE_150_io_data_2_in_bits),
    .io_data_2_out_valid(PE_150_io_data_2_out_valid),
    .io_data_2_out_bits(PE_150_io_data_2_out_bits),
    .io_data_1_in_valid(PE_150_io_data_1_in_valid),
    .io_data_1_in_bits(PE_150_io_data_1_in_bits),
    .io_data_1_out_valid(PE_150_io_data_1_out_valid),
    .io_data_1_out_bits(PE_150_io_data_1_out_bits),
    .io_data_0_in_valid(PE_150_io_data_0_in_valid),
    .io_data_0_in_bits(PE_150_io_data_0_in_bits),
    .io_data_0_out_valid(PE_150_io_data_0_out_valid),
    .io_data_0_out_bits(PE_150_io_data_0_out_bits),
    .io_sig_stat2trans(PE_150_io_sig_stat2trans)
  );
  PE PE_151 ( // @[pearray.scala 103:13]
    .clock(PE_151_clock),
    .reset(PE_151_reset),
    .io_data_2_in_valid(PE_151_io_data_2_in_valid),
    .io_data_2_in_bits(PE_151_io_data_2_in_bits),
    .io_data_2_out_valid(PE_151_io_data_2_out_valid),
    .io_data_2_out_bits(PE_151_io_data_2_out_bits),
    .io_data_1_in_valid(PE_151_io_data_1_in_valid),
    .io_data_1_in_bits(PE_151_io_data_1_in_bits),
    .io_data_1_out_valid(PE_151_io_data_1_out_valid),
    .io_data_1_out_bits(PE_151_io_data_1_out_bits),
    .io_data_0_in_valid(PE_151_io_data_0_in_valid),
    .io_data_0_in_bits(PE_151_io_data_0_in_bits),
    .io_data_0_out_valid(PE_151_io_data_0_out_valid),
    .io_data_0_out_bits(PE_151_io_data_0_out_bits),
    .io_sig_stat2trans(PE_151_io_sig_stat2trans)
  );
  PE PE_152 ( // @[pearray.scala 103:13]
    .clock(PE_152_clock),
    .reset(PE_152_reset),
    .io_data_2_in_valid(PE_152_io_data_2_in_valid),
    .io_data_2_in_bits(PE_152_io_data_2_in_bits),
    .io_data_2_out_valid(PE_152_io_data_2_out_valid),
    .io_data_2_out_bits(PE_152_io_data_2_out_bits),
    .io_data_1_in_valid(PE_152_io_data_1_in_valid),
    .io_data_1_in_bits(PE_152_io_data_1_in_bits),
    .io_data_1_out_valid(PE_152_io_data_1_out_valid),
    .io_data_1_out_bits(PE_152_io_data_1_out_bits),
    .io_data_0_in_valid(PE_152_io_data_0_in_valid),
    .io_data_0_in_bits(PE_152_io_data_0_in_bits),
    .io_data_0_out_valid(PE_152_io_data_0_out_valid),
    .io_data_0_out_bits(PE_152_io_data_0_out_bits),
    .io_sig_stat2trans(PE_152_io_sig_stat2trans)
  );
  PE PE_153 ( // @[pearray.scala 103:13]
    .clock(PE_153_clock),
    .reset(PE_153_reset),
    .io_data_2_in_valid(PE_153_io_data_2_in_valid),
    .io_data_2_in_bits(PE_153_io_data_2_in_bits),
    .io_data_2_out_valid(PE_153_io_data_2_out_valid),
    .io_data_2_out_bits(PE_153_io_data_2_out_bits),
    .io_data_1_in_valid(PE_153_io_data_1_in_valid),
    .io_data_1_in_bits(PE_153_io_data_1_in_bits),
    .io_data_1_out_valid(PE_153_io_data_1_out_valid),
    .io_data_1_out_bits(PE_153_io_data_1_out_bits),
    .io_data_0_in_valid(PE_153_io_data_0_in_valid),
    .io_data_0_in_bits(PE_153_io_data_0_in_bits),
    .io_data_0_out_valid(PE_153_io_data_0_out_valid),
    .io_data_0_out_bits(PE_153_io_data_0_out_bits),
    .io_sig_stat2trans(PE_153_io_sig_stat2trans)
  );
  PE PE_154 ( // @[pearray.scala 103:13]
    .clock(PE_154_clock),
    .reset(PE_154_reset),
    .io_data_2_in_valid(PE_154_io_data_2_in_valid),
    .io_data_2_in_bits(PE_154_io_data_2_in_bits),
    .io_data_2_out_valid(PE_154_io_data_2_out_valid),
    .io_data_2_out_bits(PE_154_io_data_2_out_bits),
    .io_data_1_in_valid(PE_154_io_data_1_in_valid),
    .io_data_1_in_bits(PE_154_io_data_1_in_bits),
    .io_data_1_out_valid(PE_154_io_data_1_out_valid),
    .io_data_1_out_bits(PE_154_io_data_1_out_bits),
    .io_data_0_in_valid(PE_154_io_data_0_in_valid),
    .io_data_0_in_bits(PE_154_io_data_0_in_bits),
    .io_data_0_out_valid(PE_154_io_data_0_out_valid),
    .io_data_0_out_bits(PE_154_io_data_0_out_bits),
    .io_sig_stat2trans(PE_154_io_sig_stat2trans)
  );
  PE PE_155 ( // @[pearray.scala 103:13]
    .clock(PE_155_clock),
    .reset(PE_155_reset),
    .io_data_2_in_valid(PE_155_io_data_2_in_valid),
    .io_data_2_in_bits(PE_155_io_data_2_in_bits),
    .io_data_2_out_valid(PE_155_io_data_2_out_valid),
    .io_data_2_out_bits(PE_155_io_data_2_out_bits),
    .io_data_1_in_valid(PE_155_io_data_1_in_valid),
    .io_data_1_in_bits(PE_155_io_data_1_in_bits),
    .io_data_1_out_valid(PE_155_io_data_1_out_valid),
    .io_data_1_out_bits(PE_155_io_data_1_out_bits),
    .io_data_0_in_valid(PE_155_io_data_0_in_valid),
    .io_data_0_in_bits(PE_155_io_data_0_in_bits),
    .io_data_0_out_valid(PE_155_io_data_0_out_valid),
    .io_data_0_out_bits(PE_155_io_data_0_out_bits),
    .io_sig_stat2trans(PE_155_io_sig_stat2trans)
  );
  PE PE_156 ( // @[pearray.scala 103:13]
    .clock(PE_156_clock),
    .reset(PE_156_reset),
    .io_data_2_in_valid(PE_156_io_data_2_in_valid),
    .io_data_2_in_bits(PE_156_io_data_2_in_bits),
    .io_data_2_out_valid(PE_156_io_data_2_out_valid),
    .io_data_2_out_bits(PE_156_io_data_2_out_bits),
    .io_data_1_in_valid(PE_156_io_data_1_in_valid),
    .io_data_1_in_bits(PE_156_io_data_1_in_bits),
    .io_data_1_out_valid(PE_156_io_data_1_out_valid),
    .io_data_1_out_bits(PE_156_io_data_1_out_bits),
    .io_data_0_in_valid(PE_156_io_data_0_in_valid),
    .io_data_0_in_bits(PE_156_io_data_0_in_bits),
    .io_data_0_out_valid(PE_156_io_data_0_out_valid),
    .io_data_0_out_bits(PE_156_io_data_0_out_bits),
    .io_sig_stat2trans(PE_156_io_sig_stat2trans)
  );
  PE PE_157 ( // @[pearray.scala 103:13]
    .clock(PE_157_clock),
    .reset(PE_157_reset),
    .io_data_2_in_valid(PE_157_io_data_2_in_valid),
    .io_data_2_in_bits(PE_157_io_data_2_in_bits),
    .io_data_2_out_valid(PE_157_io_data_2_out_valid),
    .io_data_2_out_bits(PE_157_io_data_2_out_bits),
    .io_data_1_in_valid(PE_157_io_data_1_in_valid),
    .io_data_1_in_bits(PE_157_io_data_1_in_bits),
    .io_data_1_out_valid(PE_157_io_data_1_out_valid),
    .io_data_1_out_bits(PE_157_io_data_1_out_bits),
    .io_data_0_in_valid(PE_157_io_data_0_in_valid),
    .io_data_0_in_bits(PE_157_io_data_0_in_bits),
    .io_data_0_out_valid(PE_157_io_data_0_out_valid),
    .io_data_0_out_bits(PE_157_io_data_0_out_bits),
    .io_sig_stat2trans(PE_157_io_sig_stat2trans)
  );
  PE PE_158 ( // @[pearray.scala 103:13]
    .clock(PE_158_clock),
    .reset(PE_158_reset),
    .io_data_2_in_valid(PE_158_io_data_2_in_valid),
    .io_data_2_in_bits(PE_158_io_data_2_in_bits),
    .io_data_2_out_valid(PE_158_io_data_2_out_valid),
    .io_data_2_out_bits(PE_158_io_data_2_out_bits),
    .io_data_1_in_valid(PE_158_io_data_1_in_valid),
    .io_data_1_in_bits(PE_158_io_data_1_in_bits),
    .io_data_1_out_valid(PE_158_io_data_1_out_valid),
    .io_data_1_out_bits(PE_158_io_data_1_out_bits),
    .io_data_0_in_valid(PE_158_io_data_0_in_valid),
    .io_data_0_in_bits(PE_158_io_data_0_in_bits),
    .io_data_0_out_valid(PE_158_io_data_0_out_valid),
    .io_data_0_out_bits(PE_158_io_data_0_out_bits),
    .io_sig_stat2trans(PE_158_io_sig_stat2trans)
  );
  PE PE_159 ( // @[pearray.scala 103:13]
    .clock(PE_159_clock),
    .reset(PE_159_reset),
    .io_data_2_in_valid(PE_159_io_data_2_in_valid),
    .io_data_2_in_bits(PE_159_io_data_2_in_bits),
    .io_data_2_out_valid(PE_159_io_data_2_out_valid),
    .io_data_2_out_bits(PE_159_io_data_2_out_bits),
    .io_data_1_in_valid(PE_159_io_data_1_in_valid),
    .io_data_1_in_bits(PE_159_io_data_1_in_bits),
    .io_data_1_out_valid(PE_159_io_data_1_out_valid),
    .io_data_1_out_bits(PE_159_io_data_1_out_bits),
    .io_data_0_in_valid(PE_159_io_data_0_in_valid),
    .io_data_0_in_bits(PE_159_io_data_0_in_bits),
    .io_data_0_out_valid(PE_159_io_data_0_out_valid),
    .io_data_0_out_bits(PE_159_io_data_0_out_bits),
    .io_sig_stat2trans(PE_159_io_sig_stat2trans)
  );
  PE PE_160 ( // @[pearray.scala 103:13]
    .clock(PE_160_clock),
    .reset(PE_160_reset),
    .io_data_2_in_valid(PE_160_io_data_2_in_valid),
    .io_data_2_in_bits(PE_160_io_data_2_in_bits),
    .io_data_2_out_valid(PE_160_io_data_2_out_valid),
    .io_data_2_out_bits(PE_160_io_data_2_out_bits),
    .io_data_1_in_valid(PE_160_io_data_1_in_valid),
    .io_data_1_in_bits(PE_160_io_data_1_in_bits),
    .io_data_1_out_valid(PE_160_io_data_1_out_valid),
    .io_data_1_out_bits(PE_160_io_data_1_out_bits),
    .io_data_0_in_valid(PE_160_io_data_0_in_valid),
    .io_data_0_in_bits(PE_160_io_data_0_in_bits),
    .io_data_0_out_valid(PE_160_io_data_0_out_valid),
    .io_data_0_out_bits(PE_160_io_data_0_out_bits),
    .io_sig_stat2trans(PE_160_io_sig_stat2trans)
  );
  PE PE_161 ( // @[pearray.scala 103:13]
    .clock(PE_161_clock),
    .reset(PE_161_reset),
    .io_data_2_in_valid(PE_161_io_data_2_in_valid),
    .io_data_2_in_bits(PE_161_io_data_2_in_bits),
    .io_data_2_out_valid(PE_161_io_data_2_out_valid),
    .io_data_2_out_bits(PE_161_io_data_2_out_bits),
    .io_data_1_in_valid(PE_161_io_data_1_in_valid),
    .io_data_1_in_bits(PE_161_io_data_1_in_bits),
    .io_data_1_out_valid(PE_161_io_data_1_out_valid),
    .io_data_1_out_bits(PE_161_io_data_1_out_bits),
    .io_data_0_in_valid(PE_161_io_data_0_in_valid),
    .io_data_0_in_bits(PE_161_io_data_0_in_bits),
    .io_data_0_out_valid(PE_161_io_data_0_out_valid),
    .io_data_0_out_bits(PE_161_io_data_0_out_bits),
    .io_sig_stat2trans(PE_161_io_sig_stat2trans)
  );
  PE PE_162 ( // @[pearray.scala 103:13]
    .clock(PE_162_clock),
    .reset(PE_162_reset),
    .io_data_2_in_valid(PE_162_io_data_2_in_valid),
    .io_data_2_in_bits(PE_162_io_data_2_in_bits),
    .io_data_2_out_valid(PE_162_io_data_2_out_valid),
    .io_data_2_out_bits(PE_162_io_data_2_out_bits),
    .io_data_1_in_valid(PE_162_io_data_1_in_valid),
    .io_data_1_in_bits(PE_162_io_data_1_in_bits),
    .io_data_1_out_valid(PE_162_io_data_1_out_valid),
    .io_data_1_out_bits(PE_162_io_data_1_out_bits),
    .io_data_0_in_valid(PE_162_io_data_0_in_valid),
    .io_data_0_in_bits(PE_162_io_data_0_in_bits),
    .io_data_0_out_valid(PE_162_io_data_0_out_valid),
    .io_data_0_out_bits(PE_162_io_data_0_out_bits),
    .io_sig_stat2trans(PE_162_io_sig_stat2trans)
  );
  PE PE_163 ( // @[pearray.scala 103:13]
    .clock(PE_163_clock),
    .reset(PE_163_reset),
    .io_data_2_in_valid(PE_163_io_data_2_in_valid),
    .io_data_2_in_bits(PE_163_io_data_2_in_bits),
    .io_data_2_out_valid(PE_163_io_data_2_out_valid),
    .io_data_2_out_bits(PE_163_io_data_2_out_bits),
    .io_data_1_in_valid(PE_163_io_data_1_in_valid),
    .io_data_1_in_bits(PE_163_io_data_1_in_bits),
    .io_data_1_out_valid(PE_163_io_data_1_out_valid),
    .io_data_1_out_bits(PE_163_io_data_1_out_bits),
    .io_data_0_in_valid(PE_163_io_data_0_in_valid),
    .io_data_0_in_bits(PE_163_io_data_0_in_bits),
    .io_data_0_out_valid(PE_163_io_data_0_out_valid),
    .io_data_0_out_bits(PE_163_io_data_0_out_bits),
    .io_sig_stat2trans(PE_163_io_sig_stat2trans)
  );
  PE PE_164 ( // @[pearray.scala 103:13]
    .clock(PE_164_clock),
    .reset(PE_164_reset),
    .io_data_2_in_valid(PE_164_io_data_2_in_valid),
    .io_data_2_in_bits(PE_164_io_data_2_in_bits),
    .io_data_2_out_valid(PE_164_io_data_2_out_valid),
    .io_data_2_out_bits(PE_164_io_data_2_out_bits),
    .io_data_1_in_valid(PE_164_io_data_1_in_valid),
    .io_data_1_in_bits(PE_164_io_data_1_in_bits),
    .io_data_1_out_valid(PE_164_io_data_1_out_valid),
    .io_data_1_out_bits(PE_164_io_data_1_out_bits),
    .io_data_0_in_valid(PE_164_io_data_0_in_valid),
    .io_data_0_in_bits(PE_164_io_data_0_in_bits),
    .io_data_0_out_valid(PE_164_io_data_0_out_valid),
    .io_data_0_out_bits(PE_164_io_data_0_out_bits),
    .io_sig_stat2trans(PE_164_io_sig_stat2trans)
  );
  PE PE_165 ( // @[pearray.scala 103:13]
    .clock(PE_165_clock),
    .reset(PE_165_reset),
    .io_data_2_in_valid(PE_165_io_data_2_in_valid),
    .io_data_2_in_bits(PE_165_io_data_2_in_bits),
    .io_data_2_out_valid(PE_165_io_data_2_out_valid),
    .io_data_2_out_bits(PE_165_io_data_2_out_bits),
    .io_data_1_in_valid(PE_165_io_data_1_in_valid),
    .io_data_1_in_bits(PE_165_io_data_1_in_bits),
    .io_data_1_out_valid(PE_165_io_data_1_out_valid),
    .io_data_1_out_bits(PE_165_io_data_1_out_bits),
    .io_data_0_in_valid(PE_165_io_data_0_in_valid),
    .io_data_0_in_bits(PE_165_io_data_0_in_bits),
    .io_data_0_out_valid(PE_165_io_data_0_out_valid),
    .io_data_0_out_bits(PE_165_io_data_0_out_bits),
    .io_sig_stat2trans(PE_165_io_sig_stat2trans)
  );
  PE PE_166 ( // @[pearray.scala 103:13]
    .clock(PE_166_clock),
    .reset(PE_166_reset),
    .io_data_2_in_valid(PE_166_io_data_2_in_valid),
    .io_data_2_in_bits(PE_166_io_data_2_in_bits),
    .io_data_2_out_valid(PE_166_io_data_2_out_valid),
    .io_data_2_out_bits(PE_166_io_data_2_out_bits),
    .io_data_1_in_valid(PE_166_io_data_1_in_valid),
    .io_data_1_in_bits(PE_166_io_data_1_in_bits),
    .io_data_1_out_valid(PE_166_io_data_1_out_valid),
    .io_data_1_out_bits(PE_166_io_data_1_out_bits),
    .io_data_0_in_valid(PE_166_io_data_0_in_valid),
    .io_data_0_in_bits(PE_166_io_data_0_in_bits),
    .io_data_0_out_valid(PE_166_io_data_0_out_valid),
    .io_data_0_out_bits(PE_166_io_data_0_out_bits),
    .io_sig_stat2trans(PE_166_io_sig_stat2trans)
  );
  PE PE_167 ( // @[pearray.scala 103:13]
    .clock(PE_167_clock),
    .reset(PE_167_reset),
    .io_data_2_in_valid(PE_167_io_data_2_in_valid),
    .io_data_2_in_bits(PE_167_io_data_2_in_bits),
    .io_data_2_out_valid(PE_167_io_data_2_out_valid),
    .io_data_2_out_bits(PE_167_io_data_2_out_bits),
    .io_data_1_in_valid(PE_167_io_data_1_in_valid),
    .io_data_1_in_bits(PE_167_io_data_1_in_bits),
    .io_data_1_out_valid(PE_167_io_data_1_out_valid),
    .io_data_1_out_bits(PE_167_io_data_1_out_bits),
    .io_data_0_in_valid(PE_167_io_data_0_in_valid),
    .io_data_0_in_bits(PE_167_io_data_0_in_bits),
    .io_data_0_out_valid(PE_167_io_data_0_out_valid),
    .io_data_0_out_bits(PE_167_io_data_0_out_bits),
    .io_sig_stat2trans(PE_167_io_sig_stat2trans)
  );
  PE PE_168 ( // @[pearray.scala 103:13]
    .clock(PE_168_clock),
    .reset(PE_168_reset),
    .io_data_2_in_valid(PE_168_io_data_2_in_valid),
    .io_data_2_in_bits(PE_168_io_data_2_in_bits),
    .io_data_2_out_valid(PE_168_io_data_2_out_valid),
    .io_data_2_out_bits(PE_168_io_data_2_out_bits),
    .io_data_1_in_valid(PE_168_io_data_1_in_valid),
    .io_data_1_in_bits(PE_168_io_data_1_in_bits),
    .io_data_1_out_valid(PE_168_io_data_1_out_valid),
    .io_data_1_out_bits(PE_168_io_data_1_out_bits),
    .io_data_0_in_valid(PE_168_io_data_0_in_valid),
    .io_data_0_in_bits(PE_168_io_data_0_in_bits),
    .io_data_0_out_valid(PE_168_io_data_0_out_valid),
    .io_data_0_out_bits(PE_168_io_data_0_out_bits),
    .io_sig_stat2trans(PE_168_io_sig_stat2trans)
  );
  PE PE_169 ( // @[pearray.scala 103:13]
    .clock(PE_169_clock),
    .reset(PE_169_reset),
    .io_data_2_in_valid(PE_169_io_data_2_in_valid),
    .io_data_2_in_bits(PE_169_io_data_2_in_bits),
    .io_data_2_out_valid(PE_169_io_data_2_out_valid),
    .io_data_2_out_bits(PE_169_io_data_2_out_bits),
    .io_data_1_in_valid(PE_169_io_data_1_in_valid),
    .io_data_1_in_bits(PE_169_io_data_1_in_bits),
    .io_data_1_out_valid(PE_169_io_data_1_out_valid),
    .io_data_1_out_bits(PE_169_io_data_1_out_bits),
    .io_data_0_in_valid(PE_169_io_data_0_in_valid),
    .io_data_0_in_bits(PE_169_io_data_0_in_bits),
    .io_data_0_out_valid(PE_169_io_data_0_out_valid),
    .io_data_0_out_bits(PE_169_io_data_0_out_bits),
    .io_sig_stat2trans(PE_169_io_sig_stat2trans)
  );
  PE PE_170 ( // @[pearray.scala 103:13]
    .clock(PE_170_clock),
    .reset(PE_170_reset),
    .io_data_2_in_valid(PE_170_io_data_2_in_valid),
    .io_data_2_in_bits(PE_170_io_data_2_in_bits),
    .io_data_2_out_valid(PE_170_io_data_2_out_valid),
    .io_data_2_out_bits(PE_170_io_data_2_out_bits),
    .io_data_1_in_valid(PE_170_io_data_1_in_valid),
    .io_data_1_in_bits(PE_170_io_data_1_in_bits),
    .io_data_1_out_valid(PE_170_io_data_1_out_valid),
    .io_data_1_out_bits(PE_170_io_data_1_out_bits),
    .io_data_0_in_valid(PE_170_io_data_0_in_valid),
    .io_data_0_in_bits(PE_170_io_data_0_in_bits),
    .io_data_0_out_valid(PE_170_io_data_0_out_valid),
    .io_data_0_out_bits(PE_170_io_data_0_out_bits),
    .io_sig_stat2trans(PE_170_io_sig_stat2trans)
  );
  PE PE_171 ( // @[pearray.scala 103:13]
    .clock(PE_171_clock),
    .reset(PE_171_reset),
    .io_data_2_in_valid(PE_171_io_data_2_in_valid),
    .io_data_2_in_bits(PE_171_io_data_2_in_bits),
    .io_data_2_out_valid(PE_171_io_data_2_out_valid),
    .io_data_2_out_bits(PE_171_io_data_2_out_bits),
    .io_data_1_in_valid(PE_171_io_data_1_in_valid),
    .io_data_1_in_bits(PE_171_io_data_1_in_bits),
    .io_data_1_out_valid(PE_171_io_data_1_out_valid),
    .io_data_1_out_bits(PE_171_io_data_1_out_bits),
    .io_data_0_in_valid(PE_171_io_data_0_in_valid),
    .io_data_0_in_bits(PE_171_io_data_0_in_bits),
    .io_data_0_out_valid(PE_171_io_data_0_out_valid),
    .io_data_0_out_bits(PE_171_io_data_0_out_bits),
    .io_sig_stat2trans(PE_171_io_sig_stat2trans)
  );
  PE PE_172 ( // @[pearray.scala 103:13]
    .clock(PE_172_clock),
    .reset(PE_172_reset),
    .io_data_2_in_valid(PE_172_io_data_2_in_valid),
    .io_data_2_in_bits(PE_172_io_data_2_in_bits),
    .io_data_2_out_valid(PE_172_io_data_2_out_valid),
    .io_data_2_out_bits(PE_172_io_data_2_out_bits),
    .io_data_1_in_valid(PE_172_io_data_1_in_valid),
    .io_data_1_in_bits(PE_172_io_data_1_in_bits),
    .io_data_1_out_valid(PE_172_io_data_1_out_valid),
    .io_data_1_out_bits(PE_172_io_data_1_out_bits),
    .io_data_0_in_valid(PE_172_io_data_0_in_valid),
    .io_data_0_in_bits(PE_172_io_data_0_in_bits),
    .io_data_0_out_valid(PE_172_io_data_0_out_valid),
    .io_data_0_out_bits(PE_172_io_data_0_out_bits),
    .io_sig_stat2trans(PE_172_io_sig_stat2trans)
  );
  PE PE_173 ( // @[pearray.scala 103:13]
    .clock(PE_173_clock),
    .reset(PE_173_reset),
    .io_data_2_in_valid(PE_173_io_data_2_in_valid),
    .io_data_2_in_bits(PE_173_io_data_2_in_bits),
    .io_data_2_out_valid(PE_173_io_data_2_out_valid),
    .io_data_2_out_bits(PE_173_io_data_2_out_bits),
    .io_data_1_in_valid(PE_173_io_data_1_in_valid),
    .io_data_1_in_bits(PE_173_io_data_1_in_bits),
    .io_data_1_out_valid(PE_173_io_data_1_out_valid),
    .io_data_1_out_bits(PE_173_io_data_1_out_bits),
    .io_data_0_in_valid(PE_173_io_data_0_in_valid),
    .io_data_0_in_bits(PE_173_io_data_0_in_bits),
    .io_data_0_out_valid(PE_173_io_data_0_out_valid),
    .io_data_0_out_bits(PE_173_io_data_0_out_bits),
    .io_sig_stat2trans(PE_173_io_sig_stat2trans)
  );
  PE PE_174 ( // @[pearray.scala 103:13]
    .clock(PE_174_clock),
    .reset(PE_174_reset),
    .io_data_2_in_valid(PE_174_io_data_2_in_valid),
    .io_data_2_in_bits(PE_174_io_data_2_in_bits),
    .io_data_2_out_valid(PE_174_io_data_2_out_valid),
    .io_data_2_out_bits(PE_174_io_data_2_out_bits),
    .io_data_1_in_valid(PE_174_io_data_1_in_valid),
    .io_data_1_in_bits(PE_174_io_data_1_in_bits),
    .io_data_1_out_valid(PE_174_io_data_1_out_valid),
    .io_data_1_out_bits(PE_174_io_data_1_out_bits),
    .io_data_0_in_valid(PE_174_io_data_0_in_valid),
    .io_data_0_in_bits(PE_174_io_data_0_in_bits),
    .io_data_0_out_valid(PE_174_io_data_0_out_valid),
    .io_data_0_out_bits(PE_174_io_data_0_out_bits),
    .io_sig_stat2trans(PE_174_io_sig_stat2trans)
  );
  PE PE_175 ( // @[pearray.scala 103:13]
    .clock(PE_175_clock),
    .reset(PE_175_reset),
    .io_data_2_in_valid(PE_175_io_data_2_in_valid),
    .io_data_2_in_bits(PE_175_io_data_2_in_bits),
    .io_data_2_out_valid(PE_175_io_data_2_out_valid),
    .io_data_2_out_bits(PE_175_io_data_2_out_bits),
    .io_data_1_in_valid(PE_175_io_data_1_in_valid),
    .io_data_1_in_bits(PE_175_io_data_1_in_bits),
    .io_data_1_out_valid(PE_175_io_data_1_out_valid),
    .io_data_1_out_bits(PE_175_io_data_1_out_bits),
    .io_data_0_in_valid(PE_175_io_data_0_in_valid),
    .io_data_0_in_bits(PE_175_io_data_0_in_bits),
    .io_data_0_out_valid(PE_175_io_data_0_out_valid),
    .io_data_0_out_bits(PE_175_io_data_0_out_bits),
    .io_sig_stat2trans(PE_175_io_sig_stat2trans)
  );
  PE PE_176 ( // @[pearray.scala 103:13]
    .clock(PE_176_clock),
    .reset(PE_176_reset),
    .io_data_2_in_valid(PE_176_io_data_2_in_valid),
    .io_data_2_in_bits(PE_176_io_data_2_in_bits),
    .io_data_2_out_valid(PE_176_io_data_2_out_valid),
    .io_data_2_out_bits(PE_176_io_data_2_out_bits),
    .io_data_1_in_valid(PE_176_io_data_1_in_valid),
    .io_data_1_in_bits(PE_176_io_data_1_in_bits),
    .io_data_1_out_valid(PE_176_io_data_1_out_valid),
    .io_data_1_out_bits(PE_176_io_data_1_out_bits),
    .io_data_0_in_valid(PE_176_io_data_0_in_valid),
    .io_data_0_in_bits(PE_176_io_data_0_in_bits),
    .io_data_0_out_valid(PE_176_io_data_0_out_valid),
    .io_data_0_out_bits(PE_176_io_data_0_out_bits),
    .io_sig_stat2trans(PE_176_io_sig_stat2trans)
  );
  PE PE_177 ( // @[pearray.scala 103:13]
    .clock(PE_177_clock),
    .reset(PE_177_reset),
    .io_data_2_in_valid(PE_177_io_data_2_in_valid),
    .io_data_2_in_bits(PE_177_io_data_2_in_bits),
    .io_data_2_out_valid(PE_177_io_data_2_out_valid),
    .io_data_2_out_bits(PE_177_io_data_2_out_bits),
    .io_data_1_in_valid(PE_177_io_data_1_in_valid),
    .io_data_1_in_bits(PE_177_io_data_1_in_bits),
    .io_data_1_out_valid(PE_177_io_data_1_out_valid),
    .io_data_1_out_bits(PE_177_io_data_1_out_bits),
    .io_data_0_in_valid(PE_177_io_data_0_in_valid),
    .io_data_0_in_bits(PE_177_io_data_0_in_bits),
    .io_data_0_out_valid(PE_177_io_data_0_out_valid),
    .io_data_0_out_bits(PE_177_io_data_0_out_bits),
    .io_sig_stat2trans(PE_177_io_sig_stat2trans)
  );
  PE PE_178 ( // @[pearray.scala 103:13]
    .clock(PE_178_clock),
    .reset(PE_178_reset),
    .io_data_2_in_valid(PE_178_io_data_2_in_valid),
    .io_data_2_in_bits(PE_178_io_data_2_in_bits),
    .io_data_2_out_valid(PE_178_io_data_2_out_valid),
    .io_data_2_out_bits(PE_178_io_data_2_out_bits),
    .io_data_1_in_valid(PE_178_io_data_1_in_valid),
    .io_data_1_in_bits(PE_178_io_data_1_in_bits),
    .io_data_1_out_valid(PE_178_io_data_1_out_valid),
    .io_data_1_out_bits(PE_178_io_data_1_out_bits),
    .io_data_0_in_valid(PE_178_io_data_0_in_valid),
    .io_data_0_in_bits(PE_178_io_data_0_in_bits),
    .io_data_0_out_valid(PE_178_io_data_0_out_valid),
    .io_data_0_out_bits(PE_178_io_data_0_out_bits),
    .io_sig_stat2trans(PE_178_io_sig_stat2trans)
  );
  PE PE_179 ( // @[pearray.scala 103:13]
    .clock(PE_179_clock),
    .reset(PE_179_reset),
    .io_data_2_in_valid(PE_179_io_data_2_in_valid),
    .io_data_2_in_bits(PE_179_io_data_2_in_bits),
    .io_data_2_out_valid(PE_179_io_data_2_out_valid),
    .io_data_2_out_bits(PE_179_io_data_2_out_bits),
    .io_data_1_in_valid(PE_179_io_data_1_in_valid),
    .io_data_1_in_bits(PE_179_io_data_1_in_bits),
    .io_data_1_out_valid(PE_179_io_data_1_out_valid),
    .io_data_1_out_bits(PE_179_io_data_1_out_bits),
    .io_data_0_in_valid(PE_179_io_data_0_in_valid),
    .io_data_0_in_bits(PE_179_io_data_0_in_bits),
    .io_data_0_out_valid(PE_179_io_data_0_out_valid),
    .io_data_0_out_bits(PE_179_io_data_0_out_bits),
    .io_sig_stat2trans(PE_179_io_sig_stat2trans)
  );
  PE PE_180 ( // @[pearray.scala 103:13]
    .clock(PE_180_clock),
    .reset(PE_180_reset),
    .io_data_2_in_valid(PE_180_io_data_2_in_valid),
    .io_data_2_in_bits(PE_180_io_data_2_in_bits),
    .io_data_2_out_valid(PE_180_io_data_2_out_valid),
    .io_data_2_out_bits(PE_180_io_data_2_out_bits),
    .io_data_1_in_valid(PE_180_io_data_1_in_valid),
    .io_data_1_in_bits(PE_180_io_data_1_in_bits),
    .io_data_1_out_valid(PE_180_io_data_1_out_valid),
    .io_data_1_out_bits(PE_180_io_data_1_out_bits),
    .io_data_0_in_valid(PE_180_io_data_0_in_valid),
    .io_data_0_in_bits(PE_180_io_data_0_in_bits),
    .io_data_0_out_valid(PE_180_io_data_0_out_valid),
    .io_data_0_out_bits(PE_180_io_data_0_out_bits),
    .io_sig_stat2trans(PE_180_io_sig_stat2trans)
  );
  PE PE_181 ( // @[pearray.scala 103:13]
    .clock(PE_181_clock),
    .reset(PE_181_reset),
    .io_data_2_in_valid(PE_181_io_data_2_in_valid),
    .io_data_2_in_bits(PE_181_io_data_2_in_bits),
    .io_data_2_out_valid(PE_181_io_data_2_out_valid),
    .io_data_2_out_bits(PE_181_io_data_2_out_bits),
    .io_data_1_in_valid(PE_181_io_data_1_in_valid),
    .io_data_1_in_bits(PE_181_io_data_1_in_bits),
    .io_data_1_out_valid(PE_181_io_data_1_out_valid),
    .io_data_1_out_bits(PE_181_io_data_1_out_bits),
    .io_data_0_in_valid(PE_181_io_data_0_in_valid),
    .io_data_0_in_bits(PE_181_io_data_0_in_bits),
    .io_data_0_out_valid(PE_181_io_data_0_out_valid),
    .io_data_0_out_bits(PE_181_io_data_0_out_bits),
    .io_sig_stat2trans(PE_181_io_sig_stat2trans)
  );
  PE PE_182 ( // @[pearray.scala 103:13]
    .clock(PE_182_clock),
    .reset(PE_182_reset),
    .io_data_2_in_valid(PE_182_io_data_2_in_valid),
    .io_data_2_in_bits(PE_182_io_data_2_in_bits),
    .io_data_2_out_valid(PE_182_io_data_2_out_valid),
    .io_data_2_out_bits(PE_182_io_data_2_out_bits),
    .io_data_1_in_valid(PE_182_io_data_1_in_valid),
    .io_data_1_in_bits(PE_182_io_data_1_in_bits),
    .io_data_1_out_valid(PE_182_io_data_1_out_valid),
    .io_data_1_out_bits(PE_182_io_data_1_out_bits),
    .io_data_0_in_valid(PE_182_io_data_0_in_valid),
    .io_data_0_in_bits(PE_182_io_data_0_in_bits),
    .io_data_0_out_valid(PE_182_io_data_0_out_valid),
    .io_data_0_out_bits(PE_182_io_data_0_out_bits),
    .io_sig_stat2trans(PE_182_io_sig_stat2trans)
  );
  PE PE_183 ( // @[pearray.scala 103:13]
    .clock(PE_183_clock),
    .reset(PE_183_reset),
    .io_data_2_in_valid(PE_183_io_data_2_in_valid),
    .io_data_2_in_bits(PE_183_io_data_2_in_bits),
    .io_data_2_out_valid(PE_183_io_data_2_out_valid),
    .io_data_2_out_bits(PE_183_io_data_2_out_bits),
    .io_data_1_in_valid(PE_183_io_data_1_in_valid),
    .io_data_1_in_bits(PE_183_io_data_1_in_bits),
    .io_data_1_out_valid(PE_183_io_data_1_out_valid),
    .io_data_1_out_bits(PE_183_io_data_1_out_bits),
    .io_data_0_in_valid(PE_183_io_data_0_in_valid),
    .io_data_0_in_bits(PE_183_io_data_0_in_bits),
    .io_data_0_out_valid(PE_183_io_data_0_out_valid),
    .io_data_0_out_bits(PE_183_io_data_0_out_bits),
    .io_sig_stat2trans(PE_183_io_sig_stat2trans)
  );
  PE PE_184 ( // @[pearray.scala 103:13]
    .clock(PE_184_clock),
    .reset(PE_184_reset),
    .io_data_2_in_valid(PE_184_io_data_2_in_valid),
    .io_data_2_in_bits(PE_184_io_data_2_in_bits),
    .io_data_2_out_valid(PE_184_io_data_2_out_valid),
    .io_data_2_out_bits(PE_184_io_data_2_out_bits),
    .io_data_1_in_valid(PE_184_io_data_1_in_valid),
    .io_data_1_in_bits(PE_184_io_data_1_in_bits),
    .io_data_1_out_valid(PE_184_io_data_1_out_valid),
    .io_data_1_out_bits(PE_184_io_data_1_out_bits),
    .io_data_0_in_valid(PE_184_io_data_0_in_valid),
    .io_data_0_in_bits(PE_184_io_data_0_in_bits),
    .io_data_0_out_valid(PE_184_io_data_0_out_valid),
    .io_data_0_out_bits(PE_184_io_data_0_out_bits),
    .io_sig_stat2trans(PE_184_io_sig_stat2trans)
  );
  PE PE_185 ( // @[pearray.scala 103:13]
    .clock(PE_185_clock),
    .reset(PE_185_reset),
    .io_data_2_in_valid(PE_185_io_data_2_in_valid),
    .io_data_2_in_bits(PE_185_io_data_2_in_bits),
    .io_data_2_out_valid(PE_185_io_data_2_out_valid),
    .io_data_2_out_bits(PE_185_io_data_2_out_bits),
    .io_data_1_in_valid(PE_185_io_data_1_in_valid),
    .io_data_1_in_bits(PE_185_io_data_1_in_bits),
    .io_data_1_out_valid(PE_185_io_data_1_out_valid),
    .io_data_1_out_bits(PE_185_io_data_1_out_bits),
    .io_data_0_in_valid(PE_185_io_data_0_in_valid),
    .io_data_0_in_bits(PE_185_io_data_0_in_bits),
    .io_data_0_out_valid(PE_185_io_data_0_out_valid),
    .io_data_0_out_bits(PE_185_io_data_0_out_bits),
    .io_sig_stat2trans(PE_185_io_sig_stat2trans)
  );
  PE PE_186 ( // @[pearray.scala 103:13]
    .clock(PE_186_clock),
    .reset(PE_186_reset),
    .io_data_2_in_valid(PE_186_io_data_2_in_valid),
    .io_data_2_in_bits(PE_186_io_data_2_in_bits),
    .io_data_2_out_valid(PE_186_io_data_2_out_valid),
    .io_data_2_out_bits(PE_186_io_data_2_out_bits),
    .io_data_1_in_valid(PE_186_io_data_1_in_valid),
    .io_data_1_in_bits(PE_186_io_data_1_in_bits),
    .io_data_1_out_valid(PE_186_io_data_1_out_valid),
    .io_data_1_out_bits(PE_186_io_data_1_out_bits),
    .io_data_0_in_valid(PE_186_io_data_0_in_valid),
    .io_data_0_in_bits(PE_186_io_data_0_in_bits),
    .io_data_0_out_valid(PE_186_io_data_0_out_valid),
    .io_data_0_out_bits(PE_186_io_data_0_out_bits),
    .io_sig_stat2trans(PE_186_io_sig_stat2trans)
  );
  PE PE_187 ( // @[pearray.scala 103:13]
    .clock(PE_187_clock),
    .reset(PE_187_reset),
    .io_data_2_in_valid(PE_187_io_data_2_in_valid),
    .io_data_2_in_bits(PE_187_io_data_2_in_bits),
    .io_data_2_out_valid(PE_187_io_data_2_out_valid),
    .io_data_2_out_bits(PE_187_io_data_2_out_bits),
    .io_data_1_in_valid(PE_187_io_data_1_in_valid),
    .io_data_1_in_bits(PE_187_io_data_1_in_bits),
    .io_data_1_out_valid(PE_187_io_data_1_out_valid),
    .io_data_1_out_bits(PE_187_io_data_1_out_bits),
    .io_data_0_in_valid(PE_187_io_data_0_in_valid),
    .io_data_0_in_bits(PE_187_io_data_0_in_bits),
    .io_data_0_out_valid(PE_187_io_data_0_out_valid),
    .io_data_0_out_bits(PE_187_io_data_0_out_bits),
    .io_sig_stat2trans(PE_187_io_sig_stat2trans)
  );
  PE PE_188 ( // @[pearray.scala 103:13]
    .clock(PE_188_clock),
    .reset(PE_188_reset),
    .io_data_2_in_valid(PE_188_io_data_2_in_valid),
    .io_data_2_in_bits(PE_188_io_data_2_in_bits),
    .io_data_2_out_valid(PE_188_io_data_2_out_valid),
    .io_data_2_out_bits(PE_188_io_data_2_out_bits),
    .io_data_1_in_valid(PE_188_io_data_1_in_valid),
    .io_data_1_in_bits(PE_188_io_data_1_in_bits),
    .io_data_1_out_valid(PE_188_io_data_1_out_valid),
    .io_data_1_out_bits(PE_188_io_data_1_out_bits),
    .io_data_0_in_valid(PE_188_io_data_0_in_valid),
    .io_data_0_in_bits(PE_188_io_data_0_in_bits),
    .io_data_0_out_valid(PE_188_io_data_0_out_valid),
    .io_data_0_out_bits(PE_188_io_data_0_out_bits),
    .io_sig_stat2trans(PE_188_io_sig_stat2trans)
  );
  PE PE_189 ( // @[pearray.scala 103:13]
    .clock(PE_189_clock),
    .reset(PE_189_reset),
    .io_data_2_in_valid(PE_189_io_data_2_in_valid),
    .io_data_2_in_bits(PE_189_io_data_2_in_bits),
    .io_data_2_out_valid(PE_189_io_data_2_out_valid),
    .io_data_2_out_bits(PE_189_io_data_2_out_bits),
    .io_data_1_in_valid(PE_189_io_data_1_in_valid),
    .io_data_1_in_bits(PE_189_io_data_1_in_bits),
    .io_data_1_out_valid(PE_189_io_data_1_out_valid),
    .io_data_1_out_bits(PE_189_io_data_1_out_bits),
    .io_data_0_in_valid(PE_189_io_data_0_in_valid),
    .io_data_0_in_bits(PE_189_io_data_0_in_bits),
    .io_data_0_out_valid(PE_189_io_data_0_out_valid),
    .io_data_0_out_bits(PE_189_io_data_0_out_bits),
    .io_sig_stat2trans(PE_189_io_sig_stat2trans)
  );
  PE PE_190 ( // @[pearray.scala 103:13]
    .clock(PE_190_clock),
    .reset(PE_190_reset),
    .io_data_2_in_valid(PE_190_io_data_2_in_valid),
    .io_data_2_in_bits(PE_190_io_data_2_in_bits),
    .io_data_2_out_valid(PE_190_io_data_2_out_valid),
    .io_data_2_out_bits(PE_190_io_data_2_out_bits),
    .io_data_1_in_valid(PE_190_io_data_1_in_valid),
    .io_data_1_in_bits(PE_190_io_data_1_in_bits),
    .io_data_1_out_valid(PE_190_io_data_1_out_valid),
    .io_data_1_out_bits(PE_190_io_data_1_out_bits),
    .io_data_0_in_valid(PE_190_io_data_0_in_valid),
    .io_data_0_in_bits(PE_190_io_data_0_in_bits),
    .io_data_0_out_valid(PE_190_io_data_0_out_valid),
    .io_data_0_out_bits(PE_190_io_data_0_out_bits),
    .io_sig_stat2trans(PE_190_io_sig_stat2trans)
  );
  PE PE_191 ( // @[pearray.scala 103:13]
    .clock(PE_191_clock),
    .reset(PE_191_reset),
    .io_data_2_in_valid(PE_191_io_data_2_in_valid),
    .io_data_2_in_bits(PE_191_io_data_2_in_bits),
    .io_data_2_out_valid(PE_191_io_data_2_out_valid),
    .io_data_2_out_bits(PE_191_io_data_2_out_bits),
    .io_data_1_in_valid(PE_191_io_data_1_in_valid),
    .io_data_1_in_bits(PE_191_io_data_1_in_bits),
    .io_data_1_out_valid(PE_191_io_data_1_out_valid),
    .io_data_1_out_bits(PE_191_io_data_1_out_bits),
    .io_data_0_in_valid(PE_191_io_data_0_in_valid),
    .io_data_0_in_bits(PE_191_io_data_0_in_bits),
    .io_data_0_out_valid(PE_191_io_data_0_out_valid),
    .io_data_0_out_bits(PE_191_io_data_0_out_bits),
    .io_sig_stat2trans(PE_191_io_sig_stat2trans)
  );
  PE PE_192 ( // @[pearray.scala 103:13]
    .clock(PE_192_clock),
    .reset(PE_192_reset),
    .io_data_2_in_valid(PE_192_io_data_2_in_valid),
    .io_data_2_in_bits(PE_192_io_data_2_in_bits),
    .io_data_2_out_valid(PE_192_io_data_2_out_valid),
    .io_data_2_out_bits(PE_192_io_data_2_out_bits),
    .io_data_1_in_valid(PE_192_io_data_1_in_valid),
    .io_data_1_in_bits(PE_192_io_data_1_in_bits),
    .io_data_1_out_valid(PE_192_io_data_1_out_valid),
    .io_data_1_out_bits(PE_192_io_data_1_out_bits),
    .io_data_0_in_valid(PE_192_io_data_0_in_valid),
    .io_data_0_in_bits(PE_192_io_data_0_in_bits),
    .io_data_0_out_valid(PE_192_io_data_0_out_valid),
    .io_data_0_out_bits(PE_192_io_data_0_out_bits),
    .io_sig_stat2trans(PE_192_io_sig_stat2trans)
  );
  PE PE_193 ( // @[pearray.scala 103:13]
    .clock(PE_193_clock),
    .reset(PE_193_reset),
    .io_data_2_in_valid(PE_193_io_data_2_in_valid),
    .io_data_2_in_bits(PE_193_io_data_2_in_bits),
    .io_data_2_out_valid(PE_193_io_data_2_out_valid),
    .io_data_2_out_bits(PE_193_io_data_2_out_bits),
    .io_data_1_in_valid(PE_193_io_data_1_in_valid),
    .io_data_1_in_bits(PE_193_io_data_1_in_bits),
    .io_data_1_out_valid(PE_193_io_data_1_out_valid),
    .io_data_1_out_bits(PE_193_io_data_1_out_bits),
    .io_data_0_in_valid(PE_193_io_data_0_in_valid),
    .io_data_0_in_bits(PE_193_io_data_0_in_bits),
    .io_data_0_out_valid(PE_193_io_data_0_out_valid),
    .io_data_0_out_bits(PE_193_io_data_0_out_bits),
    .io_sig_stat2trans(PE_193_io_sig_stat2trans)
  );
  PE PE_194 ( // @[pearray.scala 103:13]
    .clock(PE_194_clock),
    .reset(PE_194_reset),
    .io_data_2_in_valid(PE_194_io_data_2_in_valid),
    .io_data_2_in_bits(PE_194_io_data_2_in_bits),
    .io_data_2_out_valid(PE_194_io_data_2_out_valid),
    .io_data_2_out_bits(PE_194_io_data_2_out_bits),
    .io_data_1_in_valid(PE_194_io_data_1_in_valid),
    .io_data_1_in_bits(PE_194_io_data_1_in_bits),
    .io_data_1_out_valid(PE_194_io_data_1_out_valid),
    .io_data_1_out_bits(PE_194_io_data_1_out_bits),
    .io_data_0_in_valid(PE_194_io_data_0_in_valid),
    .io_data_0_in_bits(PE_194_io_data_0_in_bits),
    .io_data_0_out_valid(PE_194_io_data_0_out_valid),
    .io_data_0_out_bits(PE_194_io_data_0_out_bits),
    .io_sig_stat2trans(PE_194_io_sig_stat2trans)
  );
  PE PE_195 ( // @[pearray.scala 103:13]
    .clock(PE_195_clock),
    .reset(PE_195_reset),
    .io_data_2_in_valid(PE_195_io_data_2_in_valid),
    .io_data_2_in_bits(PE_195_io_data_2_in_bits),
    .io_data_2_out_valid(PE_195_io_data_2_out_valid),
    .io_data_2_out_bits(PE_195_io_data_2_out_bits),
    .io_data_1_in_valid(PE_195_io_data_1_in_valid),
    .io_data_1_in_bits(PE_195_io_data_1_in_bits),
    .io_data_1_out_valid(PE_195_io_data_1_out_valid),
    .io_data_1_out_bits(PE_195_io_data_1_out_bits),
    .io_data_0_in_valid(PE_195_io_data_0_in_valid),
    .io_data_0_in_bits(PE_195_io_data_0_in_bits),
    .io_data_0_out_valid(PE_195_io_data_0_out_valid),
    .io_data_0_out_bits(PE_195_io_data_0_out_bits),
    .io_sig_stat2trans(PE_195_io_sig_stat2trans)
  );
  PE PE_196 ( // @[pearray.scala 103:13]
    .clock(PE_196_clock),
    .reset(PE_196_reset),
    .io_data_2_in_valid(PE_196_io_data_2_in_valid),
    .io_data_2_in_bits(PE_196_io_data_2_in_bits),
    .io_data_2_out_valid(PE_196_io_data_2_out_valid),
    .io_data_2_out_bits(PE_196_io_data_2_out_bits),
    .io_data_1_in_valid(PE_196_io_data_1_in_valid),
    .io_data_1_in_bits(PE_196_io_data_1_in_bits),
    .io_data_1_out_valid(PE_196_io_data_1_out_valid),
    .io_data_1_out_bits(PE_196_io_data_1_out_bits),
    .io_data_0_in_valid(PE_196_io_data_0_in_valid),
    .io_data_0_in_bits(PE_196_io_data_0_in_bits),
    .io_data_0_out_valid(PE_196_io_data_0_out_valid),
    .io_data_0_out_bits(PE_196_io_data_0_out_bits),
    .io_sig_stat2trans(PE_196_io_sig_stat2trans)
  );
  PE PE_197 ( // @[pearray.scala 103:13]
    .clock(PE_197_clock),
    .reset(PE_197_reset),
    .io_data_2_in_valid(PE_197_io_data_2_in_valid),
    .io_data_2_in_bits(PE_197_io_data_2_in_bits),
    .io_data_2_out_valid(PE_197_io_data_2_out_valid),
    .io_data_2_out_bits(PE_197_io_data_2_out_bits),
    .io_data_1_in_valid(PE_197_io_data_1_in_valid),
    .io_data_1_in_bits(PE_197_io_data_1_in_bits),
    .io_data_1_out_valid(PE_197_io_data_1_out_valid),
    .io_data_1_out_bits(PE_197_io_data_1_out_bits),
    .io_data_0_in_valid(PE_197_io_data_0_in_valid),
    .io_data_0_in_bits(PE_197_io_data_0_in_bits),
    .io_data_0_out_valid(PE_197_io_data_0_out_valid),
    .io_data_0_out_bits(PE_197_io_data_0_out_bits),
    .io_sig_stat2trans(PE_197_io_sig_stat2trans)
  );
  PE PE_198 ( // @[pearray.scala 103:13]
    .clock(PE_198_clock),
    .reset(PE_198_reset),
    .io_data_2_in_valid(PE_198_io_data_2_in_valid),
    .io_data_2_in_bits(PE_198_io_data_2_in_bits),
    .io_data_2_out_valid(PE_198_io_data_2_out_valid),
    .io_data_2_out_bits(PE_198_io_data_2_out_bits),
    .io_data_1_in_valid(PE_198_io_data_1_in_valid),
    .io_data_1_in_bits(PE_198_io_data_1_in_bits),
    .io_data_1_out_valid(PE_198_io_data_1_out_valid),
    .io_data_1_out_bits(PE_198_io_data_1_out_bits),
    .io_data_0_in_valid(PE_198_io_data_0_in_valid),
    .io_data_0_in_bits(PE_198_io_data_0_in_bits),
    .io_data_0_out_valid(PE_198_io_data_0_out_valid),
    .io_data_0_out_bits(PE_198_io_data_0_out_bits),
    .io_sig_stat2trans(PE_198_io_sig_stat2trans)
  );
  PE PE_199 ( // @[pearray.scala 103:13]
    .clock(PE_199_clock),
    .reset(PE_199_reset),
    .io_data_2_in_valid(PE_199_io_data_2_in_valid),
    .io_data_2_in_bits(PE_199_io_data_2_in_bits),
    .io_data_2_out_valid(PE_199_io_data_2_out_valid),
    .io_data_2_out_bits(PE_199_io_data_2_out_bits),
    .io_data_1_in_valid(PE_199_io_data_1_in_valid),
    .io_data_1_in_bits(PE_199_io_data_1_in_bits),
    .io_data_1_out_valid(PE_199_io_data_1_out_valid),
    .io_data_1_out_bits(PE_199_io_data_1_out_bits),
    .io_data_0_in_valid(PE_199_io_data_0_in_valid),
    .io_data_0_in_bits(PE_199_io_data_0_in_bits),
    .io_data_0_out_valid(PE_199_io_data_0_out_valid),
    .io_data_0_out_bits(PE_199_io_data_0_out_bits),
    .io_sig_stat2trans(PE_199_io_sig_stat2trans)
  );
  PE PE_200 ( // @[pearray.scala 103:13]
    .clock(PE_200_clock),
    .reset(PE_200_reset),
    .io_data_2_in_valid(PE_200_io_data_2_in_valid),
    .io_data_2_in_bits(PE_200_io_data_2_in_bits),
    .io_data_2_out_valid(PE_200_io_data_2_out_valid),
    .io_data_2_out_bits(PE_200_io_data_2_out_bits),
    .io_data_1_in_valid(PE_200_io_data_1_in_valid),
    .io_data_1_in_bits(PE_200_io_data_1_in_bits),
    .io_data_1_out_valid(PE_200_io_data_1_out_valid),
    .io_data_1_out_bits(PE_200_io_data_1_out_bits),
    .io_data_0_in_valid(PE_200_io_data_0_in_valid),
    .io_data_0_in_bits(PE_200_io_data_0_in_bits),
    .io_data_0_out_valid(PE_200_io_data_0_out_valid),
    .io_data_0_out_bits(PE_200_io_data_0_out_bits),
    .io_sig_stat2trans(PE_200_io_sig_stat2trans)
  );
  PE PE_201 ( // @[pearray.scala 103:13]
    .clock(PE_201_clock),
    .reset(PE_201_reset),
    .io_data_2_in_valid(PE_201_io_data_2_in_valid),
    .io_data_2_in_bits(PE_201_io_data_2_in_bits),
    .io_data_2_out_valid(PE_201_io_data_2_out_valid),
    .io_data_2_out_bits(PE_201_io_data_2_out_bits),
    .io_data_1_in_valid(PE_201_io_data_1_in_valid),
    .io_data_1_in_bits(PE_201_io_data_1_in_bits),
    .io_data_1_out_valid(PE_201_io_data_1_out_valid),
    .io_data_1_out_bits(PE_201_io_data_1_out_bits),
    .io_data_0_in_valid(PE_201_io_data_0_in_valid),
    .io_data_0_in_bits(PE_201_io_data_0_in_bits),
    .io_data_0_out_valid(PE_201_io_data_0_out_valid),
    .io_data_0_out_bits(PE_201_io_data_0_out_bits),
    .io_sig_stat2trans(PE_201_io_sig_stat2trans)
  );
  PE PE_202 ( // @[pearray.scala 103:13]
    .clock(PE_202_clock),
    .reset(PE_202_reset),
    .io_data_2_in_valid(PE_202_io_data_2_in_valid),
    .io_data_2_in_bits(PE_202_io_data_2_in_bits),
    .io_data_2_out_valid(PE_202_io_data_2_out_valid),
    .io_data_2_out_bits(PE_202_io_data_2_out_bits),
    .io_data_1_in_valid(PE_202_io_data_1_in_valid),
    .io_data_1_in_bits(PE_202_io_data_1_in_bits),
    .io_data_1_out_valid(PE_202_io_data_1_out_valid),
    .io_data_1_out_bits(PE_202_io_data_1_out_bits),
    .io_data_0_in_valid(PE_202_io_data_0_in_valid),
    .io_data_0_in_bits(PE_202_io_data_0_in_bits),
    .io_data_0_out_valid(PE_202_io_data_0_out_valid),
    .io_data_0_out_bits(PE_202_io_data_0_out_bits),
    .io_sig_stat2trans(PE_202_io_sig_stat2trans)
  );
  PE PE_203 ( // @[pearray.scala 103:13]
    .clock(PE_203_clock),
    .reset(PE_203_reset),
    .io_data_2_in_valid(PE_203_io_data_2_in_valid),
    .io_data_2_in_bits(PE_203_io_data_2_in_bits),
    .io_data_2_out_valid(PE_203_io_data_2_out_valid),
    .io_data_2_out_bits(PE_203_io_data_2_out_bits),
    .io_data_1_in_valid(PE_203_io_data_1_in_valid),
    .io_data_1_in_bits(PE_203_io_data_1_in_bits),
    .io_data_1_out_valid(PE_203_io_data_1_out_valid),
    .io_data_1_out_bits(PE_203_io_data_1_out_bits),
    .io_data_0_in_valid(PE_203_io_data_0_in_valid),
    .io_data_0_in_bits(PE_203_io_data_0_in_bits),
    .io_data_0_out_valid(PE_203_io_data_0_out_valid),
    .io_data_0_out_bits(PE_203_io_data_0_out_bits),
    .io_sig_stat2trans(PE_203_io_sig_stat2trans)
  );
  PE PE_204 ( // @[pearray.scala 103:13]
    .clock(PE_204_clock),
    .reset(PE_204_reset),
    .io_data_2_in_valid(PE_204_io_data_2_in_valid),
    .io_data_2_in_bits(PE_204_io_data_2_in_bits),
    .io_data_2_out_valid(PE_204_io_data_2_out_valid),
    .io_data_2_out_bits(PE_204_io_data_2_out_bits),
    .io_data_1_in_valid(PE_204_io_data_1_in_valid),
    .io_data_1_in_bits(PE_204_io_data_1_in_bits),
    .io_data_1_out_valid(PE_204_io_data_1_out_valid),
    .io_data_1_out_bits(PE_204_io_data_1_out_bits),
    .io_data_0_in_valid(PE_204_io_data_0_in_valid),
    .io_data_0_in_bits(PE_204_io_data_0_in_bits),
    .io_data_0_out_valid(PE_204_io_data_0_out_valid),
    .io_data_0_out_bits(PE_204_io_data_0_out_bits),
    .io_sig_stat2trans(PE_204_io_sig_stat2trans)
  );
  PE PE_205 ( // @[pearray.scala 103:13]
    .clock(PE_205_clock),
    .reset(PE_205_reset),
    .io_data_2_in_valid(PE_205_io_data_2_in_valid),
    .io_data_2_in_bits(PE_205_io_data_2_in_bits),
    .io_data_2_out_valid(PE_205_io_data_2_out_valid),
    .io_data_2_out_bits(PE_205_io_data_2_out_bits),
    .io_data_1_in_valid(PE_205_io_data_1_in_valid),
    .io_data_1_in_bits(PE_205_io_data_1_in_bits),
    .io_data_1_out_valid(PE_205_io_data_1_out_valid),
    .io_data_1_out_bits(PE_205_io_data_1_out_bits),
    .io_data_0_in_valid(PE_205_io_data_0_in_valid),
    .io_data_0_in_bits(PE_205_io_data_0_in_bits),
    .io_data_0_out_valid(PE_205_io_data_0_out_valid),
    .io_data_0_out_bits(PE_205_io_data_0_out_bits),
    .io_sig_stat2trans(PE_205_io_sig_stat2trans)
  );
  PE PE_206 ( // @[pearray.scala 103:13]
    .clock(PE_206_clock),
    .reset(PE_206_reset),
    .io_data_2_in_valid(PE_206_io_data_2_in_valid),
    .io_data_2_in_bits(PE_206_io_data_2_in_bits),
    .io_data_2_out_valid(PE_206_io_data_2_out_valid),
    .io_data_2_out_bits(PE_206_io_data_2_out_bits),
    .io_data_1_in_valid(PE_206_io_data_1_in_valid),
    .io_data_1_in_bits(PE_206_io_data_1_in_bits),
    .io_data_1_out_valid(PE_206_io_data_1_out_valid),
    .io_data_1_out_bits(PE_206_io_data_1_out_bits),
    .io_data_0_in_valid(PE_206_io_data_0_in_valid),
    .io_data_0_in_bits(PE_206_io_data_0_in_bits),
    .io_data_0_out_valid(PE_206_io_data_0_out_valid),
    .io_data_0_out_bits(PE_206_io_data_0_out_bits),
    .io_sig_stat2trans(PE_206_io_sig_stat2trans)
  );
  PE PE_207 ( // @[pearray.scala 103:13]
    .clock(PE_207_clock),
    .reset(PE_207_reset),
    .io_data_2_in_valid(PE_207_io_data_2_in_valid),
    .io_data_2_in_bits(PE_207_io_data_2_in_bits),
    .io_data_2_out_valid(PE_207_io_data_2_out_valid),
    .io_data_2_out_bits(PE_207_io_data_2_out_bits),
    .io_data_1_in_valid(PE_207_io_data_1_in_valid),
    .io_data_1_in_bits(PE_207_io_data_1_in_bits),
    .io_data_1_out_valid(PE_207_io_data_1_out_valid),
    .io_data_1_out_bits(PE_207_io_data_1_out_bits),
    .io_data_0_in_valid(PE_207_io_data_0_in_valid),
    .io_data_0_in_bits(PE_207_io_data_0_in_bits),
    .io_data_0_out_valid(PE_207_io_data_0_out_valid),
    .io_data_0_out_bits(PE_207_io_data_0_out_bits),
    .io_sig_stat2trans(PE_207_io_sig_stat2trans)
  );
  PE PE_208 ( // @[pearray.scala 103:13]
    .clock(PE_208_clock),
    .reset(PE_208_reset),
    .io_data_2_in_valid(PE_208_io_data_2_in_valid),
    .io_data_2_in_bits(PE_208_io_data_2_in_bits),
    .io_data_2_out_valid(PE_208_io_data_2_out_valid),
    .io_data_2_out_bits(PE_208_io_data_2_out_bits),
    .io_data_1_in_valid(PE_208_io_data_1_in_valid),
    .io_data_1_in_bits(PE_208_io_data_1_in_bits),
    .io_data_1_out_valid(PE_208_io_data_1_out_valid),
    .io_data_1_out_bits(PE_208_io_data_1_out_bits),
    .io_data_0_in_valid(PE_208_io_data_0_in_valid),
    .io_data_0_in_bits(PE_208_io_data_0_in_bits),
    .io_data_0_out_valid(PE_208_io_data_0_out_valid),
    .io_data_0_out_bits(PE_208_io_data_0_out_bits),
    .io_sig_stat2trans(PE_208_io_sig_stat2trans)
  );
  PE PE_209 ( // @[pearray.scala 103:13]
    .clock(PE_209_clock),
    .reset(PE_209_reset),
    .io_data_2_in_valid(PE_209_io_data_2_in_valid),
    .io_data_2_in_bits(PE_209_io_data_2_in_bits),
    .io_data_2_out_valid(PE_209_io_data_2_out_valid),
    .io_data_2_out_bits(PE_209_io_data_2_out_bits),
    .io_data_1_in_valid(PE_209_io_data_1_in_valid),
    .io_data_1_in_bits(PE_209_io_data_1_in_bits),
    .io_data_1_out_valid(PE_209_io_data_1_out_valid),
    .io_data_1_out_bits(PE_209_io_data_1_out_bits),
    .io_data_0_in_valid(PE_209_io_data_0_in_valid),
    .io_data_0_in_bits(PE_209_io_data_0_in_bits),
    .io_data_0_out_valid(PE_209_io_data_0_out_valid),
    .io_data_0_out_bits(PE_209_io_data_0_out_bits),
    .io_sig_stat2trans(PE_209_io_sig_stat2trans)
  );
  PE PE_210 ( // @[pearray.scala 103:13]
    .clock(PE_210_clock),
    .reset(PE_210_reset),
    .io_data_2_in_valid(PE_210_io_data_2_in_valid),
    .io_data_2_in_bits(PE_210_io_data_2_in_bits),
    .io_data_2_out_valid(PE_210_io_data_2_out_valid),
    .io_data_2_out_bits(PE_210_io_data_2_out_bits),
    .io_data_1_in_valid(PE_210_io_data_1_in_valid),
    .io_data_1_in_bits(PE_210_io_data_1_in_bits),
    .io_data_1_out_valid(PE_210_io_data_1_out_valid),
    .io_data_1_out_bits(PE_210_io_data_1_out_bits),
    .io_data_0_in_valid(PE_210_io_data_0_in_valid),
    .io_data_0_in_bits(PE_210_io_data_0_in_bits),
    .io_data_0_out_valid(PE_210_io_data_0_out_valid),
    .io_data_0_out_bits(PE_210_io_data_0_out_bits),
    .io_sig_stat2trans(PE_210_io_sig_stat2trans)
  );
  PE PE_211 ( // @[pearray.scala 103:13]
    .clock(PE_211_clock),
    .reset(PE_211_reset),
    .io_data_2_in_valid(PE_211_io_data_2_in_valid),
    .io_data_2_in_bits(PE_211_io_data_2_in_bits),
    .io_data_2_out_valid(PE_211_io_data_2_out_valid),
    .io_data_2_out_bits(PE_211_io_data_2_out_bits),
    .io_data_1_in_valid(PE_211_io_data_1_in_valid),
    .io_data_1_in_bits(PE_211_io_data_1_in_bits),
    .io_data_1_out_valid(PE_211_io_data_1_out_valid),
    .io_data_1_out_bits(PE_211_io_data_1_out_bits),
    .io_data_0_in_valid(PE_211_io_data_0_in_valid),
    .io_data_0_in_bits(PE_211_io_data_0_in_bits),
    .io_data_0_out_valid(PE_211_io_data_0_out_valid),
    .io_data_0_out_bits(PE_211_io_data_0_out_bits),
    .io_sig_stat2trans(PE_211_io_sig_stat2trans)
  );
  PE PE_212 ( // @[pearray.scala 103:13]
    .clock(PE_212_clock),
    .reset(PE_212_reset),
    .io_data_2_in_valid(PE_212_io_data_2_in_valid),
    .io_data_2_in_bits(PE_212_io_data_2_in_bits),
    .io_data_2_out_valid(PE_212_io_data_2_out_valid),
    .io_data_2_out_bits(PE_212_io_data_2_out_bits),
    .io_data_1_in_valid(PE_212_io_data_1_in_valid),
    .io_data_1_in_bits(PE_212_io_data_1_in_bits),
    .io_data_1_out_valid(PE_212_io_data_1_out_valid),
    .io_data_1_out_bits(PE_212_io_data_1_out_bits),
    .io_data_0_in_valid(PE_212_io_data_0_in_valid),
    .io_data_0_in_bits(PE_212_io_data_0_in_bits),
    .io_data_0_out_valid(PE_212_io_data_0_out_valid),
    .io_data_0_out_bits(PE_212_io_data_0_out_bits),
    .io_sig_stat2trans(PE_212_io_sig_stat2trans)
  );
  PE PE_213 ( // @[pearray.scala 103:13]
    .clock(PE_213_clock),
    .reset(PE_213_reset),
    .io_data_2_in_valid(PE_213_io_data_2_in_valid),
    .io_data_2_in_bits(PE_213_io_data_2_in_bits),
    .io_data_2_out_valid(PE_213_io_data_2_out_valid),
    .io_data_2_out_bits(PE_213_io_data_2_out_bits),
    .io_data_1_in_valid(PE_213_io_data_1_in_valid),
    .io_data_1_in_bits(PE_213_io_data_1_in_bits),
    .io_data_1_out_valid(PE_213_io_data_1_out_valid),
    .io_data_1_out_bits(PE_213_io_data_1_out_bits),
    .io_data_0_in_valid(PE_213_io_data_0_in_valid),
    .io_data_0_in_bits(PE_213_io_data_0_in_bits),
    .io_data_0_out_valid(PE_213_io_data_0_out_valid),
    .io_data_0_out_bits(PE_213_io_data_0_out_bits),
    .io_sig_stat2trans(PE_213_io_sig_stat2trans)
  );
  PE PE_214 ( // @[pearray.scala 103:13]
    .clock(PE_214_clock),
    .reset(PE_214_reset),
    .io_data_2_in_valid(PE_214_io_data_2_in_valid),
    .io_data_2_in_bits(PE_214_io_data_2_in_bits),
    .io_data_2_out_valid(PE_214_io_data_2_out_valid),
    .io_data_2_out_bits(PE_214_io_data_2_out_bits),
    .io_data_1_in_valid(PE_214_io_data_1_in_valid),
    .io_data_1_in_bits(PE_214_io_data_1_in_bits),
    .io_data_1_out_valid(PE_214_io_data_1_out_valid),
    .io_data_1_out_bits(PE_214_io_data_1_out_bits),
    .io_data_0_in_valid(PE_214_io_data_0_in_valid),
    .io_data_0_in_bits(PE_214_io_data_0_in_bits),
    .io_data_0_out_valid(PE_214_io_data_0_out_valid),
    .io_data_0_out_bits(PE_214_io_data_0_out_bits),
    .io_sig_stat2trans(PE_214_io_sig_stat2trans)
  );
  PE PE_215 ( // @[pearray.scala 103:13]
    .clock(PE_215_clock),
    .reset(PE_215_reset),
    .io_data_2_in_valid(PE_215_io_data_2_in_valid),
    .io_data_2_in_bits(PE_215_io_data_2_in_bits),
    .io_data_2_out_valid(PE_215_io_data_2_out_valid),
    .io_data_2_out_bits(PE_215_io_data_2_out_bits),
    .io_data_1_in_valid(PE_215_io_data_1_in_valid),
    .io_data_1_in_bits(PE_215_io_data_1_in_bits),
    .io_data_1_out_valid(PE_215_io_data_1_out_valid),
    .io_data_1_out_bits(PE_215_io_data_1_out_bits),
    .io_data_0_in_valid(PE_215_io_data_0_in_valid),
    .io_data_0_in_bits(PE_215_io_data_0_in_bits),
    .io_data_0_out_valid(PE_215_io_data_0_out_valid),
    .io_data_0_out_bits(PE_215_io_data_0_out_bits),
    .io_sig_stat2trans(PE_215_io_sig_stat2trans)
  );
  PE PE_216 ( // @[pearray.scala 103:13]
    .clock(PE_216_clock),
    .reset(PE_216_reset),
    .io_data_2_in_valid(PE_216_io_data_2_in_valid),
    .io_data_2_in_bits(PE_216_io_data_2_in_bits),
    .io_data_2_out_valid(PE_216_io_data_2_out_valid),
    .io_data_2_out_bits(PE_216_io_data_2_out_bits),
    .io_data_1_in_valid(PE_216_io_data_1_in_valid),
    .io_data_1_in_bits(PE_216_io_data_1_in_bits),
    .io_data_1_out_valid(PE_216_io_data_1_out_valid),
    .io_data_1_out_bits(PE_216_io_data_1_out_bits),
    .io_data_0_in_valid(PE_216_io_data_0_in_valid),
    .io_data_0_in_bits(PE_216_io_data_0_in_bits),
    .io_data_0_out_valid(PE_216_io_data_0_out_valid),
    .io_data_0_out_bits(PE_216_io_data_0_out_bits),
    .io_sig_stat2trans(PE_216_io_sig_stat2trans)
  );
  PE PE_217 ( // @[pearray.scala 103:13]
    .clock(PE_217_clock),
    .reset(PE_217_reset),
    .io_data_2_in_valid(PE_217_io_data_2_in_valid),
    .io_data_2_in_bits(PE_217_io_data_2_in_bits),
    .io_data_2_out_valid(PE_217_io_data_2_out_valid),
    .io_data_2_out_bits(PE_217_io_data_2_out_bits),
    .io_data_1_in_valid(PE_217_io_data_1_in_valid),
    .io_data_1_in_bits(PE_217_io_data_1_in_bits),
    .io_data_1_out_valid(PE_217_io_data_1_out_valid),
    .io_data_1_out_bits(PE_217_io_data_1_out_bits),
    .io_data_0_in_valid(PE_217_io_data_0_in_valid),
    .io_data_0_in_bits(PE_217_io_data_0_in_bits),
    .io_data_0_out_valid(PE_217_io_data_0_out_valid),
    .io_data_0_out_bits(PE_217_io_data_0_out_bits),
    .io_sig_stat2trans(PE_217_io_sig_stat2trans)
  );
  PE PE_218 ( // @[pearray.scala 103:13]
    .clock(PE_218_clock),
    .reset(PE_218_reset),
    .io_data_2_in_valid(PE_218_io_data_2_in_valid),
    .io_data_2_in_bits(PE_218_io_data_2_in_bits),
    .io_data_2_out_valid(PE_218_io_data_2_out_valid),
    .io_data_2_out_bits(PE_218_io_data_2_out_bits),
    .io_data_1_in_valid(PE_218_io_data_1_in_valid),
    .io_data_1_in_bits(PE_218_io_data_1_in_bits),
    .io_data_1_out_valid(PE_218_io_data_1_out_valid),
    .io_data_1_out_bits(PE_218_io_data_1_out_bits),
    .io_data_0_in_valid(PE_218_io_data_0_in_valid),
    .io_data_0_in_bits(PE_218_io_data_0_in_bits),
    .io_data_0_out_valid(PE_218_io_data_0_out_valid),
    .io_data_0_out_bits(PE_218_io_data_0_out_bits),
    .io_sig_stat2trans(PE_218_io_sig_stat2trans)
  );
  PE PE_219 ( // @[pearray.scala 103:13]
    .clock(PE_219_clock),
    .reset(PE_219_reset),
    .io_data_2_in_valid(PE_219_io_data_2_in_valid),
    .io_data_2_in_bits(PE_219_io_data_2_in_bits),
    .io_data_2_out_valid(PE_219_io_data_2_out_valid),
    .io_data_2_out_bits(PE_219_io_data_2_out_bits),
    .io_data_1_in_valid(PE_219_io_data_1_in_valid),
    .io_data_1_in_bits(PE_219_io_data_1_in_bits),
    .io_data_1_out_valid(PE_219_io_data_1_out_valid),
    .io_data_1_out_bits(PE_219_io_data_1_out_bits),
    .io_data_0_in_valid(PE_219_io_data_0_in_valid),
    .io_data_0_in_bits(PE_219_io_data_0_in_bits),
    .io_data_0_out_valid(PE_219_io_data_0_out_valid),
    .io_data_0_out_bits(PE_219_io_data_0_out_bits),
    .io_sig_stat2trans(PE_219_io_sig_stat2trans)
  );
  PE PE_220 ( // @[pearray.scala 103:13]
    .clock(PE_220_clock),
    .reset(PE_220_reset),
    .io_data_2_in_valid(PE_220_io_data_2_in_valid),
    .io_data_2_in_bits(PE_220_io_data_2_in_bits),
    .io_data_2_out_valid(PE_220_io_data_2_out_valid),
    .io_data_2_out_bits(PE_220_io_data_2_out_bits),
    .io_data_1_in_valid(PE_220_io_data_1_in_valid),
    .io_data_1_in_bits(PE_220_io_data_1_in_bits),
    .io_data_1_out_valid(PE_220_io_data_1_out_valid),
    .io_data_1_out_bits(PE_220_io_data_1_out_bits),
    .io_data_0_in_valid(PE_220_io_data_0_in_valid),
    .io_data_0_in_bits(PE_220_io_data_0_in_bits),
    .io_data_0_out_valid(PE_220_io_data_0_out_valid),
    .io_data_0_out_bits(PE_220_io_data_0_out_bits),
    .io_sig_stat2trans(PE_220_io_sig_stat2trans)
  );
  PE PE_221 ( // @[pearray.scala 103:13]
    .clock(PE_221_clock),
    .reset(PE_221_reset),
    .io_data_2_in_valid(PE_221_io_data_2_in_valid),
    .io_data_2_in_bits(PE_221_io_data_2_in_bits),
    .io_data_2_out_valid(PE_221_io_data_2_out_valid),
    .io_data_2_out_bits(PE_221_io_data_2_out_bits),
    .io_data_1_in_valid(PE_221_io_data_1_in_valid),
    .io_data_1_in_bits(PE_221_io_data_1_in_bits),
    .io_data_1_out_valid(PE_221_io_data_1_out_valid),
    .io_data_1_out_bits(PE_221_io_data_1_out_bits),
    .io_data_0_in_valid(PE_221_io_data_0_in_valid),
    .io_data_0_in_bits(PE_221_io_data_0_in_bits),
    .io_data_0_out_valid(PE_221_io_data_0_out_valid),
    .io_data_0_out_bits(PE_221_io_data_0_out_bits),
    .io_sig_stat2trans(PE_221_io_sig_stat2trans)
  );
  PE PE_222 ( // @[pearray.scala 103:13]
    .clock(PE_222_clock),
    .reset(PE_222_reset),
    .io_data_2_in_valid(PE_222_io_data_2_in_valid),
    .io_data_2_in_bits(PE_222_io_data_2_in_bits),
    .io_data_2_out_valid(PE_222_io_data_2_out_valid),
    .io_data_2_out_bits(PE_222_io_data_2_out_bits),
    .io_data_1_in_valid(PE_222_io_data_1_in_valid),
    .io_data_1_in_bits(PE_222_io_data_1_in_bits),
    .io_data_1_out_valid(PE_222_io_data_1_out_valid),
    .io_data_1_out_bits(PE_222_io_data_1_out_bits),
    .io_data_0_in_valid(PE_222_io_data_0_in_valid),
    .io_data_0_in_bits(PE_222_io_data_0_in_bits),
    .io_data_0_out_valid(PE_222_io_data_0_out_valid),
    .io_data_0_out_bits(PE_222_io_data_0_out_bits),
    .io_sig_stat2trans(PE_222_io_sig_stat2trans)
  );
  PE PE_223 ( // @[pearray.scala 103:13]
    .clock(PE_223_clock),
    .reset(PE_223_reset),
    .io_data_2_in_valid(PE_223_io_data_2_in_valid),
    .io_data_2_in_bits(PE_223_io_data_2_in_bits),
    .io_data_2_out_valid(PE_223_io_data_2_out_valid),
    .io_data_2_out_bits(PE_223_io_data_2_out_bits),
    .io_data_1_in_valid(PE_223_io_data_1_in_valid),
    .io_data_1_in_bits(PE_223_io_data_1_in_bits),
    .io_data_1_out_valid(PE_223_io_data_1_out_valid),
    .io_data_1_out_bits(PE_223_io_data_1_out_bits),
    .io_data_0_in_valid(PE_223_io_data_0_in_valid),
    .io_data_0_in_bits(PE_223_io_data_0_in_bits),
    .io_data_0_out_valid(PE_223_io_data_0_out_valid),
    .io_data_0_out_bits(PE_223_io_data_0_out_bits),
    .io_sig_stat2trans(PE_223_io_sig_stat2trans)
  );
  PE PE_224 ( // @[pearray.scala 103:13]
    .clock(PE_224_clock),
    .reset(PE_224_reset),
    .io_data_2_in_valid(PE_224_io_data_2_in_valid),
    .io_data_2_in_bits(PE_224_io_data_2_in_bits),
    .io_data_2_out_valid(PE_224_io_data_2_out_valid),
    .io_data_2_out_bits(PE_224_io_data_2_out_bits),
    .io_data_1_in_valid(PE_224_io_data_1_in_valid),
    .io_data_1_in_bits(PE_224_io_data_1_in_bits),
    .io_data_1_out_valid(PE_224_io_data_1_out_valid),
    .io_data_1_out_bits(PE_224_io_data_1_out_bits),
    .io_data_0_in_valid(PE_224_io_data_0_in_valid),
    .io_data_0_in_bits(PE_224_io_data_0_in_bits),
    .io_data_0_out_valid(PE_224_io_data_0_out_valid),
    .io_data_0_out_bits(PE_224_io_data_0_out_bits),
    .io_sig_stat2trans(PE_224_io_sig_stat2trans)
  );
  PE PE_225 ( // @[pearray.scala 103:13]
    .clock(PE_225_clock),
    .reset(PE_225_reset),
    .io_data_2_in_valid(PE_225_io_data_2_in_valid),
    .io_data_2_in_bits(PE_225_io_data_2_in_bits),
    .io_data_2_out_valid(PE_225_io_data_2_out_valid),
    .io_data_2_out_bits(PE_225_io_data_2_out_bits),
    .io_data_1_in_valid(PE_225_io_data_1_in_valid),
    .io_data_1_in_bits(PE_225_io_data_1_in_bits),
    .io_data_1_out_valid(PE_225_io_data_1_out_valid),
    .io_data_1_out_bits(PE_225_io_data_1_out_bits),
    .io_data_0_in_valid(PE_225_io_data_0_in_valid),
    .io_data_0_in_bits(PE_225_io_data_0_in_bits),
    .io_data_0_out_valid(PE_225_io_data_0_out_valid),
    .io_data_0_out_bits(PE_225_io_data_0_out_bits),
    .io_sig_stat2trans(PE_225_io_sig_stat2trans)
  );
  PE PE_226 ( // @[pearray.scala 103:13]
    .clock(PE_226_clock),
    .reset(PE_226_reset),
    .io_data_2_in_valid(PE_226_io_data_2_in_valid),
    .io_data_2_in_bits(PE_226_io_data_2_in_bits),
    .io_data_2_out_valid(PE_226_io_data_2_out_valid),
    .io_data_2_out_bits(PE_226_io_data_2_out_bits),
    .io_data_1_in_valid(PE_226_io_data_1_in_valid),
    .io_data_1_in_bits(PE_226_io_data_1_in_bits),
    .io_data_1_out_valid(PE_226_io_data_1_out_valid),
    .io_data_1_out_bits(PE_226_io_data_1_out_bits),
    .io_data_0_in_valid(PE_226_io_data_0_in_valid),
    .io_data_0_in_bits(PE_226_io_data_0_in_bits),
    .io_data_0_out_valid(PE_226_io_data_0_out_valid),
    .io_data_0_out_bits(PE_226_io_data_0_out_bits),
    .io_sig_stat2trans(PE_226_io_sig_stat2trans)
  );
  PE PE_227 ( // @[pearray.scala 103:13]
    .clock(PE_227_clock),
    .reset(PE_227_reset),
    .io_data_2_in_valid(PE_227_io_data_2_in_valid),
    .io_data_2_in_bits(PE_227_io_data_2_in_bits),
    .io_data_2_out_valid(PE_227_io_data_2_out_valid),
    .io_data_2_out_bits(PE_227_io_data_2_out_bits),
    .io_data_1_in_valid(PE_227_io_data_1_in_valid),
    .io_data_1_in_bits(PE_227_io_data_1_in_bits),
    .io_data_1_out_valid(PE_227_io_data_1_out_valid),
    .io_data_1_out_bits(PE_227_io_data_1_out_bits),
    .io_data_0_in_valid(PE_227_io_data_0_in_valid),
    .io_data_0_in_bits(PE_227_io_data_0_in_bits),
    .io_data_0_out_valid(PE_227_io_data_0_out_valid),
    .io_data_0_out_bits(PE_227_io_data_0_out_bits),
    .io_sig_stat2trans(PE_227_io_sig_stat2trans)
  );
  PE PE_228 ( // @[pearray.scala 103:13]
    .clock(PE_228_clock),
    .reset(PE_228_reset),
    .io_data_2_in_valid(PE_228_io_data_2_in_valid),
    .io_data_2_in_bits(PE_228_io_data_2_in_bits),
    .io_data_2_out_valid(PE_228_io_data_2_out_valid),
    .io_data_2_out_bits(PE_228_io_data_2_out_bits),
    .io_data_1_in_valid(PE_228_io_data_1_in_valid),
    .io_data_1_in_bits(PE_228_io_data_1_in_bits),
    .io_data_1_out_valid(PE_228_io_data_1_out_valid),
    .io_data_1_out_bits(PE_228_io_data_1_out_bits),
    .io_data_0_in_valid(PE_228_io_data_0_in_valid),
    .io_data_0_in_bits(PE_228_io_data_0_in_bits),
    .io_data_0_out_valid(PE_228_io_data_0_out_valid),
    .io_data_0_out_bits(PE_228_io_data_0_out_bits),
    .io_sig_stat2trans(PE_228_io_sig_stat2trans)
  );
  PE PE_229 ( // @[pearray.scala 103:13]
    .clock(PE_229_clock),
    .reset(PE_229_reset),
    .io_data_2_in_valid(PE_229_io_data_2_in_valid),
    .io_data_2_in_bits(PE_229_io_data_2_in_bits),
    .io_data_2_out_valid(PE_229_io_data_2_out_valid),
    .io_data_2_out_bits(PE_229_io_data_2_out_bits),
    .io_data_1_in_valid(PE_229_io_data_1_in_valid),
    .io_data_1_in_bits(PE_229_io_data_1_in_bits),
    .io_data_1_out_valid(PE_229_io_data_1_out_valid),
    .io_data_1_out_bits(PE_229_io_data_1_out_bits),
    .io_data_0_in_valid(PE_229_io_data_0_in_valid),
    .io_data_0_in_bits(PE_229_io_data_0_in_bits),
    .io_data_0_out_valid(PE_229_io_data_0_out_valid),
    .io_data_0_out_bits(PE_229_io_data_0_out_bits),
    .io_sig_stat2trans(PE_229_io_sig_stat2trans)
  );
  PE PE_230 ( // @[pearray.scala 103:13]
    .clock(PE_230_clock),
    .reset(PE_230_reset),
    .io_data_2_in_valid(PE_230_io_data_2_in_valid),
    .io_data_2_in_bits(PE_230_io_data_2_in_bits),
    .io_data_2_out_valid(PE_230_io_data_2_out_valid),
    .io_data_2_out_bits(PE_230_io_data_2_out_bits),
    .io_data_1_in_valid(PE_230_io_data_1_in_valid),
    .io_data_1_in_bits(PE_230_io_data_1_in_bits),
    .io_data_1_out_valid(PE_230_io_data_1_out_valid),
    .io_data_1_out_bits(PE_230_io_data_1_out_bits),
    .io_data_0_in_valid(PE_230_io_data_0_in_valid),
    .io_data_0_in_bits(PE_230_io_data_0_in_bits),
    .io_data_0_out_valid(PE_230_io_data_0_out_valid),
    .io_data_0_out_bits(PE_230_io_data_0_out_bits),
    .io_sig_stat2trans(PE_230_io_sig_stat2trans)
  );
  PE PE_231 ( // @[pearray.scala 103:13]
    .clock(PE_231_clock),
    .reset(PE_231_reset),
    .io_data_2_in_valid(PE_231_io_data_2_in_valid),
    .io_data_2_in_bits(PE_231_io_data_2_in_bits),
    .io_data_2_out_valid(PE_231_io_data_2_out_valid),
    .io_data_2_out_bits(PE_231_io_data_2_out_bits),
    .io_data_1_in_valid(PE_231_io_data_1_in_valid),
    .io_data_1_in_bits(PE_231_io_data_1_in_bits),
    .io_data_1_out_valid(PE_231_io_data_1_out_valid),
    .io_data_1_out_bits(PE_231_io_data_1_out_bits),
    .io_data_0_in_valid(PE_231_io_data_0_in_valid),
    .io_data_0_in_bits(PE_231_io_data_0_in_bits),
    .io_data_0_out_valid(PE_231_io_data_0_out_valid),
    .io_data_0_out_bits(PE_231_io_data_0_out_bits),
    .io_sig_stat2trans(PE_231_io_sig_stat2trans)
  );
  PE PE_232 ( // @[pearray.scala 103:13]
    .clock(PE_232_clock),
    .reset(PE_232_reset),
    .io_data_2_in_valid(PE_232_io_data_2_in_valid),
    .io_data_2_in_bits(PE_232_io_data_2_in_bits),
    .io_data_2_out_valid(PE_232_io_data_2_out_valid),
    .io_data_2_out_bits(PE_232_io_data_2_out_bits),
    .io_data_1_in_valid(PE_232_io_data_1_in_valid),
    .io_data_1_in_bits(PE_232_io_data_1_in_bits),
    .io_data_1_out_valid(PE_232_io_data_1_out_valid),
    .io_data_1_out_bits(PE_232_io_data_1_out_bits),
    .io_data_0_in_valid(PE_232_io_data_0_in_valid),
    .io_data_0_in_bits(PE_232_io_data_0_in_bits),
    .io_data_0_out_valid(PE_232_io_data_0_out_valid),
    .io_data_0_out_bits(PE_232_io_data_0_out_bits),
    .io_sig_stat2trans(PE_232_io_sig_stat2trans)
  );
  PE PE_233 ( // @[pearray.scala 103:13]
    .clock(PE_233_clock),
    .reset(PE_233_reset),
    .io_data_2_in_valid(PE_233_io_data_2_in_valid),
    .io_data_2_in_bits(PE_233_io_data_2_in_bits),
    .io_data_2_out_valid(PE_233_io_data_2_out_valid),
    .io_data_2_out_bits(PE_233_io_data_2_out_bits),
    .io_data_1_in_valid(PE_233_io_data_1_in_valid),
    .io_data_1_in_bits(PE_233_io_data_1_in_bits),
    .io_data_1_out_valid(PE_233_io_data_1_out_valid),
    .io_data_1_out_bits(PE_233_io_data_1_out_bits),
    .io_data_0_in_valid(PE_233_io_data_0_in_valid),
    .io_data_0_in_bits(PE_233_io_data_0_in_bits),
    .io_data_0_out_valid(PE_233_io_data_0_out_valid),
    .io_data_0_out_bits(PE_233_io_data_0_out_bits),
    .io_sig_stat2trans(PE_233_io_sig_stat2trans)
  );
  PE PE_234 ( // @[pearray.scala 103:13]
    .clock(PE_234_clock),
    .reset(PE_234_reset),
    .io_data_2_in_valid(PE_234_io_data_2_in_valid),
    .io_data_2_in_bits(PE_234_io_data_2_in_bits),
    .io_data_2_out_valid(PE_234_io_data_2_out_valid),
    .io_data_2_out_bits(PE_234_io_data_2_out_bits),
    .io_data_1_in_valid(PE_234_io_data_1_in_valid),
    .io_data_1_in_bits(PE_234_io_data_1_in_bits),
    .io_data_1_out_valid(PE_234_io_data_1_out_valid),
    .io_data_1_out_bits(PE_234_io_data_1_out_bits),
    .io_data_0_in_valid(PE_234_io_data_0_in_valid),
    .io_data_0_in_bits(PE_234_io_data_0_in_bits),
    .io_data_0_out_valid(PE_234_io_data_0_out_valid),
    .io_data_0_out_bits(PE_234_io_data_0_out_bits),
    .io_sig_stat2trans(PE_234_io_sig_stat2trans)
  );
  PE PE_235 ( // @[pearray.scala 103:13]
    .clock(PE_235_clock),
    .reset(PE_235_reset),
    .io_data_2_in_valid(PE_235_io_data_2_in_valid),
    .io_data_2_in_bits(PE_235_io_data_2_in_bits),
    .io_data_2_out_valid(PE_235_io_data_2_out_valid),
    .io_data_2_out_bits(PE_235_io_data_2_out_bits),
    .io_data_1_in_valid(PE_235_io_data_1_in_valid),
    .io_data_1_in_bits(PE_235_io_data_1_in_bits),
    .io_data_1_out_valid(PE_235_io_data_1_out_valid),
    .io_data_1_out_bits(PE_235_io_data_1_out_bits),
    .io_data_0_in_valid(PE_235_io_data_0_in_valid),
    .io_data_0_in_bits(PE_235_io_data_0_in_bits),
    .io_data_0_out_valid(PE_235_io_data_0_out_valid),
    .io_data_0_out_bits(PE_235_io_data_0_out_bits),
    .io_sig_stat2trans(PE_235_io_sig_stat2trans)
  );
  PE PE_236 ( // @[pearray.scala 103:13]
    .clock(PE_236_clock),
    .reset(PE_236_reset),
    .io_data_2_in_valid(PE_236_io_data_2_in_valid),
    .io_data_2_in_bits(PE_236_io_data_2_in_bits),
    .io_data_2_out_valid(PE_236_io_data_2_out_valid),
    .io_data_2_out_bits(PE_236_io_data_2_out_bits),
    .io_data_1_in_valid(PE_236_io_data_1_in_valid),
    .io_data_1_in_bits(PE_236_io_data_1_in_bits),
    .io_data_1_out_valid(PE_236_io_data_1_out_valid),
    .io_data_1_out_bits(PE_236_io_data_1_out_bits),
    .io_data_0_in_valid(PE_236_io_data_0_in_valid),
    .io_data_0_in_bits(PE_236_io_data_0_in_bits),
    .io_data_0_out_valid(PE_236_io_data_0_out_valid),
    .io_data_0_out_bits(PE_236_io_data_0_out_bits),
    .io_sig_stat2trans(PE_236_io_sig_stat2trans)
  );
  PE PE_237 ( // @[pearray.scala 103:13]
    .clock(PE_237_clock),
    .reset(PE_237_reset),
    .io_data_2_in_valid(PE_237_io_data_2_in_valid),
    .io_data_2_in_bits(PE_237_io_data_2_in_bits),
    .io_data_2_out_valid(PE_237_io_data_2_out_valid),
    .io_data_2_out_bits(PE_237_io_data_2_out_bits),
    .io_data_1_in_valid(PE_237_io_data_1_in_valid),
    .io_data_1_in_bits(PE_237_io_data_1_in_bits),
    .io_data_1_out_valid(PE_237_io_data_1_out_valid),
    .io_data_1_out_bits(PE_237_io_data_1_out_bits),
    .io_data_0_in_valid(PE_237_io_data_0_in_valid),
    .io_data_0_in_bits(PE_237_io_data_0_in_bits),
    .io_data_0_out_valid(PE_237_io_data_0_out_valid),
    .io_data_0_out_bits(PE_237_io_data_0_out_bits),
    .io_sig_stat2trans(PE_237_io_sig_stat2trans)
  );
  PE PE_238 ( // @[pearray.scala 103:13]
    .clock(PE_238_clock),
    .reset(PE_238_reset),
    .io_data_2_in_valid(PE_238_io_data_2_in_valid),
    .io_data_2_in_bits(PE_238_io_data_2_in_bits),
    .io_data_2_out_valid(PE_238_io_data_2_out_valid),
    .io_data_2_out_bits(PE_238_io_data_2_out_bits),
    .io_data_1_in_valid(PE_238_io_data_1_in_valid),
    .io_data_1_in_bits(PE_238_io_data_1_in_bits),
    .io_data_1_out_valid(PE_238_io_data_1_out_valid),
    .io_data_1_out_bits(PE_238_io_data_1_out_bits),
    .io_data_0_in_valid(PE_238_io_data_0_in_valid),
    .io_data_0_in_bits(PE_238_io_data_0_in_bits),
    .io_data_0_out_valid(PE_238_io_data_0_out_valid),
    .io_data_0_out_bits(PE_238_io_data_0_out_bits),
    .io_sig_stat2trans(PE_238_io_sig_stat2trans)
  );
  PE PE_239 ( // @[pearray.scala 103:13]
    .clock(PE_239_clock),
    .reset(PE_239_reset),
    .io_data_2_in_valid(PE_239_io_data_2_in_valid),
    .io_data_2_in_bits(PE_239_io_data_2_in_bits),
    .io_data_2_out_valid(PE_239_io_data_2_out_valid),
    .io_data_2_out_bits(PE_239_io_data_2_out_bits),
    .io_data_1_in_valid(PE_239_io_data_1_in_valid),
    .io_data_1_in_bits(PE_239_io_data_1_in_bits),
    .io_data_1_out_valid(PE_239_io_data_1_out_valid),
    .io_data_1_out_bits(PE_239_io_data_1_out_bits),
    .io_data_0_in_valid(PE_239_io_data_0_in_valid),
    .io_data_0_in_bits(PE_239_io_data_0_in_bits),
    .io_data_0_out_valid(PE_239_io_data_0_out_valid),
    .io_data_0_out_bits(PE_239_io_data_0_out_bits),
    .io_sig_stat2trans(PE_239_io_sig_stat2trans)
  );
  PE PE_240 ( // @[pearray.scala 103:13]
    .clock(PE_240_clock),
    .reset(PE_240_reset),
    .io_data_2_in_valid(PE_240_io_data_2_in_valid),
    .io_data_2_in_bits(PE_240_io_data_2_in_bits),
    .io_data_2_out_valid(PE_240_io_data_2_out_valid),
    .io_data_2_out_bits(PE_240_io_data_2_out_bits),
    .io_data_1_in_valid(PE_240_io_data_1_in_valid),
    .io_data_1_in_bits(PE_240_io_data_1_in_bits),
    .io_data_1_out_valid(PE_240_io_data_1_out_valid),
    .io_data_1_out_bits(PE_240_io_data_1_out_bits),
    .io_data_0_in_valid(PE_240_io_data_0_in_valid),
    .io_data_0_in_bits(PE_240_io_data_0_in_bits),
    .io_data_0_out_valid(PE_240_io_data_0_out_valid),
    .io_data_0_out_bits(PE_240_io_data_0_out_bits),
    .io_sig_stat2trans(PE_240_io_sig_stat2trans)
  );
  PE PE_241 ( // @[pearray.scala 103:13]
    .clock(PE_241_clock),
    .reset(PE_241_reset),
    .io_data_2_in_valid(PE_241_io_data_2_in_valid),
    .io_data_2_in_bits(PE_241_io_data_2_in_bits),
    .io_data_2_out_valid(PE_241_io_data_2_out_valid),
    .io_data_2_out_bits(PE_241_io_data_2_out_bits),
    .io_data_1_in_valid(PE_241_io_data_1_in_valid),
    .io_data_1_in_bits(PE_241_io_data_1_in_bits),
    .io_data_1_out_valid(PE_241_io_data_1_out_valid),
    .io_data_1_out_bits(PE_241_io_data_1_out_bits),
    .io_data_0_in_valid(PE_241_io_data_0_in_valid),
    .io_data_0_in_bits(PE_241_io_data_0_in_bits),
    .io_data_0_out_valid(PE_241_io_data_0_out_valid),
    .io_data_0_out_bits(PE_241_io_data_0_out_bits),
    .io_sig_stat2trans(PE_241_io_sig_stat2trans)
  );
  PE PE_242 ( // @[pearray.scala 103:13]
    .clock(PE_242_clock),
    .reset(PE_242_reset),
    .io_data_2_in_valid(PE_242_io_data_2_in_valid),
    .io_data_2_in_bits(PE_242_io_data_2_in_bits),
    .io_data_2_out_valid(PE_242_io_data_2_out_valid),
    .io_data_2_out_bits(PE_242_io_data_2_out_bits),
    .io_data_1_in_valid(PE_242_io_data_1_in_valid),
    .io_data_1_in_bits(PE_242_io_data_1_in_bits),
    .io_data_1_out_valid(PE_242_io_data_1_out_valid),
    .io_data_1_out_bits(PE_242_io_data_1_out_bits),
    .io_data_0_in_valid(PE_242_io_data_0_in_valid),
    .io_data_0_in_bits(PE_242_io_data_0_in_bits),
    .io_data_0_out_valid(PE_242_io_data_0_out_valid),
    .io_data_0_out_bits(PE_242_io_data_0_out_bits),
    .io_sig_stat2trans(PE_242_io_sig_stat2trans)
  );
  PE PE_243 ( // @[pearray.scala 103:13]
    .clock(PE_243_clock),
    .reset(PE_243_reset),
    .io_data_2_in_valid(PE_243_io_data_2_in_valid),
    .io_data_2_in_bits(PE_243_io_data_2_in_bits),
    .io_data_2_out_valid(PE_243_io_data_2_out_valid),
    .io_data_2_out_bits(PE_243_io_data_2_out_bits),
    .io_data_1_in_valid(PE_243_io_data_1_in_valid),
    .io_data_1_in_bits(PE_243_io_data_1_in_bits),
    .io_data_1_out_valid(PE_243_io_data_1_out_valid),
    .io_data_1_out_bits(PE_243_io_data_1_out_bits),
    .io_data_0_in_valid(PE_243_io_data_0_in_valid),
    .io_data_0_in_bits(PE_243_io_data_0_in_bits),
    .io_data_0_out_valid(PE_243_io_data_0_out_valid),
    .io_data_0_out_bits(PE_243_io_data_0_out_bits),
    .io_sig_stat2trans(PE_243_io_sig_stat2trans)
  );
  PE PE_244 ( // @[pearray.scala 103:13]
    .clock(PE_244_clock),
    .reset(PE_244_reset),
    .io_data_2_in_valid(PE_244_io_data_2_in_valid),
    .io_data_2_in_bits(PE_244_io_data_2_in_bits),
    .io_data_2_out_valid(PE_244_io_data_2_out_valid),
    .io_data_2_out_bits(PE_244_io_data_2_out_bits),
    .io_data_1_in_valid(PE_244_io_data_1_in_valid),
    .io_data_1_in_bits(PE_244_io_data_1_in_bits),
    .io_data_1_out_valid(PE_244_io_data_1_out_valid),
    .io_data_1_out_bits(PE_244_io_data_1_out_bits),
    .io_data_0_in_valid(PE_244_io_data_0_in_valid),
    .io_data_0_in_bits(PE_244_io_data_0_in_bits),
    .io_data_0_out_valid(PE_244_io_data_0_out_valid),
    .io_data_0_out_bits(PE_244_io_data_0_out_bits),
    .io_sig_stat2trans(PE_244_io_sig_stat2trans)
  );
  PE PE_245 ( // @[pearray.scala 103:13]
    .clock(PE_245_clock),
    .reset(PE_245_reset),
    .io_data_2_in_valid(PE_245_io_data_2_in_valid),
    .io_data_2_in_bits(PE_245_io_data_2_in_bits),
    .io_data_2_out_valid(PE_245_io_data_2_out_valid),
    .io_data_2_out_bits(PE_245_io_data_2_out_bits),
    .io_data_1_in_valid(PE_245_io_data_1_in_valid),
    .io_data_1_in_bits(PE_245_io_data_1_in_bits),
    .io_data_1_out_valid(PE_245_io_data_1_out_valid),
    .io_data_1_out_bits(PE_245_io_data_1_out_bits),
    .io_data_0_in_valid(PE_245_io_data_0_in_valid),
    .io_data_0_in_bits(PE_245_io_data_0_in_bits),
    .io_data_0_out_valid(PE_245_io_data_0_out_valid),
    .io_data_0_out_bits(PE_245_io_data_0_out_bits),
    .io_sig_stat2trans(PE_245_io_sig_stat2trans)
  );
  PE PE_246 ( // @[pearray.scala 103:13]
    .clock(PE_246_clock),
    .reset(PE_246_reset),
    .io_data_2_in_valid(PE_246_io_data_2_in_valid),
    .io_data_2_in_bits(PE_246_io_data_2_in_bits),
    .io_data_2_out_valid(PE_246_io_data_2_out_valid),
    .io_data_2_out_bits(PE_246_io_data_2_out_bits),
    .io_data_1_in_valid(PE_246_io_data_1_in_valid),
    .io_data_1_in_bits(PE_246_io_data_1_in_bits),
    .io_data_1_out_valid(PE_246_io_data_1_out_valid),
    .io_data_1_out_bits(PE_246_io_data_1_out_bits),
    .io_data_0_in_valid(PE_246_io_data_0_in_valid),
    .io_data_0_in_bits(PE_246_io_data_0_in_bits),
    .io_data_0_out_valid(PE_246_io_data_0_out_valid),
    .io_data_0_out_bits(PE_246_io_data_0_out_bits),
    .io_sig_stat2trans(PE_246_io_sig_stat2trans)
  );
  PE PE_247 ( // @[pearray.scala 103:13]
    .clock(PE_247_clock),
    .reset(PE_247_reset),
    .io_data_2_in_valid(PE_247_io_data_2_in_valid),
    .io_data_2_in_bits(PE_247_io_data_2_in_bits),
    .io_data_2_out_valid(PE_247_io_data_2_out_valid),
    .io_data_2_out_bits(PE_247_io_data_2_out_bits),
    .io_data_1_in_valid(PE_247_io_data_1_in_valid),
    .io_data_1_in_bits(PE_247_io_data_1_in_bits),
    .io_data_1_out_valid(PE_247_io_data_1_out_valid),
    .io_data_1_out_bits(PE_247_io_data_1_out_bits),
    .io_data_0_in_valid(PE_247_io_data_0_in_valid),
    .io_data_0_in_bits(PE_247_io_data_0_in_bits),
    .io_data_0_out_valid(PE_247_io_data_0_out_valid),
    .io_data_0_out_bits(PE_247_io_data_0_out_bits),
    .io_sig_stat2trans(PE_247_io_sig_stat2trans)
  );
  PE PE_248 ( // @[pearray.scala 103:13]
    .clock(PE_248_clock),
    .reset(PE_248_reset),
    .io_data_2_in_valid(PE_248_io_data_2_in_valid),
    .io_data_2_in_bits(PE_248_io_data_2_in_bits),
    .io_data_2_out_valid(PE_248_io_data_2_out_valid),
    .io_data_2_out_bits(PE_248_io_data_2_out_bits),
    .io_data_1_in_valid(PE_248_io_data_1_in_valid),
    .io_data_1_in_bits(PE_248_io_data_1_in_bits),
    .io_data_1_out_valid(PE_248_io_data_1_out_valid),
    .io_data_1_out_bits(PE_248_io_data_1_out_bits),
    .io_data_0_in_valid(PE_248_io_data_0_in_valid),
    .io_data_0_in_bits(PE_248_io_data_0_in_bits),
    .io_data_0_out_valid(PE_248_io_data_0_out_valid),
    .io_data_0_out_bits(PE_248_io_data_0_out_bits),
    .io_sig_stat2trans(PE_248_io_sig_stat2trans)
  );
  PE PE_249 ( // @[pearray.scala 103:13]
    .clock(PE_249_clock),
    .reset(PE_249_reset),
    .io_data_2_in_valid(PE_249_io_data_2_in_valid),
    .io_data_2_in_bits(PE_249_io_data_2_in_bits),
    .io_data_2_out_valid(PE_249_io_data_2_out_valid),
    .io_data_2_out_bits(PE_249_io_data_2_out_bits),
    .io_data_1_in_valid(PE_249_io_data_1_in_valid),
    .io_data_1_in_bits(PE_249_io_data_1_in_bits),
    .io_data_1_out_valid(PE_249_io_data_1_out_valid),
    .io_data_1_out_bits(PE_249_io_data_1_out_bits),
    .io_data_0_in_valid(PE_249_io_data_0_in_valid),
    .io_data_0_in_bits(PE_249_io_data_0_in_bits),
    .io_data_0_out_valid(PE_249_io_data_0_out_valid),
    .io_data_0_out_bits(PE_249_io_data_0_out_bits),
    .io_sig_stat2trans(PE_249_io_sig_stat2trans)
  );
  PE PE_250 ( // @[pearray.scala 103:13]
    .clock(PE_250_clock),
    .reset(PE_250_reset),
    .io_data_2_in_valid(PE_250_io_data_2_in_valid),
    .io_data_2_in_bits(PE_250_io_data_2_in_bits),
    .io_data_2_out_valid(PE_250_io_data_2_out_valid),
    .io_data_2_out_bits(PE_250_io_data_2_out_bits),
    .io_data_1_in_valid(PE_250_io_data_1_in_valid),
    .io_data_1_in_bits(PE_250_io_data_1_in_bits),
    .io_data_1_out_valid(PE_250_io_data_1_out_valid),
    .io_data_1_out_bits(PE_250_io_data_1_out_bits),
    .io_data_0_in_valid(PE_250_io_data_0_in_valid),
    .io_data_0_in_bits(PE_250_io_data_0_in_bits),
    .io_data_0_out_valid(PE_250_io_data_0_out_valid),
    .io_data_0_out_bits(PE_250_io_data_0_out_bits),
    .io_sig_stat2trans(PE_250_io_sig_stat2trans)
  );
  PE PE_251 ( // @[pearray.scala 103:13]
    .clock(PE_251_clock),
    .reset(PE_251_reset),
    .io_data_2_in_valid(PE_251_io_data_2_in_valid),
    .io_data_2_in_bits(PE_251_io_data_2_in_bits),
    .io_data_2_out_valid(PE_251_io_data_2_out_valid),
    .io_data_2_out_bits(PE_251_io_data_2_out_bits),
    .io_data_1_in_valid(PE_251_io_data_1_in_valid),
    .io_data_1_in_bits(PE_251_io_data_1_in_bits),
    .io_data_1_out_valid(PE_251_io_data_1_out_valid),
    .io_data_1_out_bits(PE_251_io_data_1_out_bits),
    .io_data_0_in_valid(PE_251_io_data_0_in_valid),
    .io_data_0_in_bits(PE_251_io_data_0_in_bits),
    .io_data_0_out_valid(PE_251_io_data_0_out_valid),
    .io_data_0_out_bits(PE_251_io_data_0_out_bits),
    .io_sig_stat2trans(PE_251_io_sig_stat2trans)
  );
  PE PE_252 ( // @[pearray.scala 103:13]
    .clock(PE_252_clock),
    .reset(PE_252_reset),
    .io_data_2_in_valid(PE_252_io_data_2_in_valid),
    .io_data_2_in_bits(PE_252_io_data_2_in_bits),
    .io_data_2_out_valid(PE_252_io_data_2_out_valid),
    .io_data_2_out_bits(PE_252_io_data_2_out_bits),
    .io_data_1_in_valid(PE_252_io_data_1_in_valid),
    .io_data_1_in_bits(PE_252_io_data_1_in_bits),
    .io_data_1_out_valid(PE_252_io_data_1_out_valid),
    .io_data_1_out_bits(PE_252_io_data_1_out_bits),
    .io_data_0_in_valid(PE_252_io_data_0_in_valid),
    .io_data_0_in_bits(PE_252_io_data_0_in_bits),
    .io_data_0_out_valid(PE_252_io_data_0_out_valid),
    .io_data_0_out_bits(PE_252_io_data_0_out_bits),
    .io_sig_stat2trans(PE_252_io_sig_stat2trans)
  );
  PE PE_253 ( // @[pearray.scala 103:13]
    .clock(PE_253_clock),
    .reset(PE_253_reset),
    .io_data_2_in_valid(PE_253_io_data_2_in_valid),
    .io_data_2_in_bits(PE_253_io_data_2_in_bits),
    .io_data_2_out_valid(PE_253_io_data_2_out_valid),
    .io_data_2_out_bits(PE_253_io_data_2_out_bits),
    .io_data_1_in_valid(PE_253_io_data_1_in_valid),
    .io_data_1_in_bits(PE_253_io_data_1_in_bits),
    .io_data_1_out_valid(PE_253_io_data_1_out_valid),
    .io_data_1_out_bits(PE_253_io_data_1_out_bits),
    .io_data_0_in_valid(PE_253_io_data_0_in_valid),
    .io_data_0_in_bits(PE_253_io_data_0_in_bits),
    .io_data_0_out_valid(PE_253_io_data_0_out_valid),
    .io_data_0_out_bits(PE_253_io_data_0_out_bits),
    .io_sig_stat2trans(PE_253_io_sig_stat2trans)
  );
  PE PE_254 ( // @[pearray.scala 103:13]
    .clock(PE_254_clock),
    .reset(PE_254_reset),
    .io_data_2_in_valid(PE_254_io_data_2_in_valid),
    .io_data_2_in_bits(PE_254_io_data_2_in_bits),
    .io_data_2_out_valid(PE_254_io_data_2_out_valid),
    .io_data_2_out_bits(PE_254_io_data_2_out_bits),
    .io_data_1_in_valid(PE_254_io_data_1_in_valid),
    .io_data_1_in_bits(PE_254_io_data_1_in_bits),
    .io_data_1_out_valid(PE_254_io_data_1_out_valid),
    .io_data_1_out_bits(PE_254_io_data_1_out_bits),
    .io_data_0_in_valid(PE_254_io_data_0_in_valid),
    .io_data_0_in_bits(PE_254_io_data_0_in_bits),
    .io_data_0_out_valid(PE_254_io_data_0_out_valid),
    .io_data_0_out_bits(PE_254_io_data_0_out_bits),
    .io_sig_stat2trans(PE_254_io_sig_stat2trans)
  );
  PE PE_255 ( // @[pearray.scala 103:13]
    .clock(PE_255_clock),
    .reset(PE_255_reset),
    .io_data_2_in_valid(PE_255_io_data_2_in_valid),
    .io_data_2_in_bits(PE_255_io_data_2_in_bits),
    .io_data_2_out_valid(PE_255_io_data_2_out_valid),
    .io_data_2_out_bits(PE_255_io_data_2_out_bits),
    .io_data_1_in_valid(PE_255_io_data_1_in_valid),
    .io_data_1_in_bits(PE_255_io_data_1_in_bits),
    .io_data_1_out_valid(PE_255_io_data_1_out_valid),
    .io_data_1_out_bits(PE_255_io_data_1_out_bits),
    .io_data_0_in_valid(PE_255_io_data_0_in_valid),
    .io_data_0_in_bits(PE_255_io_data_0_in_bits),
    .io_data_0_out_valid(PE_255_io_data_0_out_valid),
    .io_data_0_out_bits(PE_255_io_data_0_out_bits),
    .io_sig_stat2trans(PE_255_io_sig_stat2trans)
  );
  PENetwork PENetwork ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_io_to_mem_bits)
  );
  PENetwork PENetwork_1 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_1_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_1_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_1_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_1_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_1_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_1_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_1_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_1_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_1_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_1_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_1_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_1_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_1_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_1_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_1_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_1_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_1_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_1_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_1_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_1_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_1_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_1_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_1_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_1_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_1_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_1_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_1_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_1_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_1_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_1_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_1_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_1_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_1_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_1_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_1_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_1_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_1_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_1_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_1_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_1_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_1_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_1_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_1_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_1_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_1_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_1_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_1_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_1_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_1_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_1_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_1_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_1_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_1_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_1_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_1_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_1_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_1_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_1_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_1_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_1_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_1_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_1_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_1_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_1_io_to_mem_bits)
  );
  PENetwork PENetwork_2 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_2_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_2_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_2_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_2_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_2_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_2_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_2_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_2_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_2_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_2_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_2_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_2_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_2_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_2_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_2_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_2_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_2_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_2_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_2_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_2_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_2_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_2_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_2_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_2_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_2_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_2_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_2_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_2_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_2_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_2_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_2_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_2_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_2_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_2_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_2_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_2_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_2_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_2_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_2_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_2_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_2_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_2_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_2_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_2_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_2_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_2_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_2_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_2_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_2_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_2_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_2_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_2_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_2_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_2_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_2_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_2_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_2_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_2_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_2_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_2_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_2_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_2_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_2_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_2_io_to_mem_bits)
  );
  PENetwork PENetwork_3 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_3_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_3_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_3_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_3_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_3_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_3_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_3_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_3_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_3_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_3_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_3_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_3_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_3_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_3_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_3_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_3_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_3_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_3_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_3_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_3_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_3_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_3_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_3_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_3_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_3_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_3_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_3_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_3_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_3_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_3_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_3_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_3_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_3_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_3_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_3_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_3_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_3_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_3_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_3_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_3_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_3_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_3_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_3_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_3_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_3_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_3_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_3_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_3_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_3_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_3_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_3_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_3_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_3_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_3_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_3_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_3_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_3_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_3_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_3_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_3_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_3_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_3_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_3_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_3_io_to_mem_bits)
  );
  PENetwork PENetwork_4 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_4_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_4_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_4_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_4_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_4_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_4_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_4_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_4_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_4_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_4_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_4_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_4_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_4_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_4_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_4_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_4_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_4_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_4_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_4_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_4_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_4_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_4_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_4_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_4_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_4_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_4_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_4_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_4_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_4_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_4_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_4_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_4_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_4_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_4_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_4_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_4_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_4_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_4_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_4_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_4_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_4_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_4_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_4_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_4_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_4_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_4_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_4_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_4_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_4_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_4_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_4_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_4_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_4_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_4_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_4_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_4_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_4_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_4_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_4_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_4_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_4_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_4_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_4_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_4_io_to_mem_bits)
  );
  PENetwork PENetwork_5 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_5_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_5_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_5_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_5_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_5_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_5_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_5_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_5_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_5_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_5_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_5_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_5_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_5_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_5_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_5_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_5_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_5_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_5_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_5_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_5_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_5_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_5_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_5_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_5_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_5_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_5_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_5_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_5_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_5_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_5_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_5_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_5_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_5_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_5_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_5_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_5_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_5_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_5_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_5_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_5_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_5_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_5_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_5_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_5_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_5_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_5_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_5_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_5_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_5_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_5_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_5_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_5_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_5_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_5_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_5_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_5_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_5_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_5_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_5_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_5_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_5_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_5_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_5_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_5_io_to_mem_bits)
  );
  PENetwork PENetwork_6 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_6_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_6_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_6_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_6_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_6_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_6_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_6_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_6_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_6_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_6_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_6_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_6_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_6_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_6_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_6_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_6_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_6_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_6_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_6_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_6_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_6_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_6_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_6_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_6_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_6_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_6_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_6_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_6_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_6_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_6_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_6_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_6_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_6_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_6_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_6_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_6_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_6_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_6_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_6_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_6_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_6_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_6_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_6_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_6_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_6_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_6_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_6_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_6_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_6_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_6_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_6_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_6_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_6_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_6_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_6_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_6_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_6_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_6_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_6_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_6_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_6_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_6_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_6_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_6_io_to_mem_bits)
  );
  PENetwork PENetwork_7 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_7_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_7_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_7_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_7_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_7_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_7_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_7_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_7_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_7_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_7_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_7_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_7_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_7_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_7_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_7_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_7_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_7_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_7_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_7_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_7_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_7_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_7_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_7_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_7_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_7_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_7_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_7_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_7_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_7_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_7_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_7_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_7_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_7_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_7_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_7_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_7_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_7_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_7_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_7_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_7_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_7_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_7_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_7_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_7_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_7_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_7_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_7_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_7_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_7_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_7_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_7_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_7_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_7_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_7_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_7_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_7_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_7_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_7_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_7_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_7_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_7_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_7_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_7_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_7_io_to_mem_bits)
  );
  PENetwork PENetwork_8 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_8_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_8_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_8_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_8_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_8_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_8_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_8_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_8_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_8_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_8_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_8_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_8_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_8_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_8_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_8_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_8_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_8_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_8_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_8_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_8_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_8_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_8_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_8_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_8_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_8_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_8_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_8_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_8_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_8_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_8_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_8_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_8_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_8_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_8_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_8_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_8_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_8_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_8_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_8_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_8_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_8_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_8_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_8_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_8_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_8_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_8_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_8_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_8_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_8_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_8_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_8_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_8_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_8_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_8_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_8_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_8_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_8_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_8_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_8_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_8_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_8_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_8_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_8_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_8_io_to_mem_bits)
  );
  PENetwork PENetwork_9 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_9_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_9_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_9_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_9_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_9_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_9_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_9_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_9_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_9_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_9_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_9_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_9_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_9_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_9_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_9_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_9_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_9_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_9_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_9_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_9_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_9_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_9_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_9_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_9_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_9_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_9_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_9_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_9_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_9_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_9_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_9_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_9_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_9_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_9_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_9_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_9_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_9_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_9_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_9_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_9_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_9_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_9_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_9_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_9_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_9_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_9_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_9_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_9_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_9_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_9_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_9_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_9_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_9_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_9_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_9_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_9_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_9_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_9_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_9_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_9_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_9_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_9_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_9_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_9_io_to_mem_bits)
  );
  PENetwork PENetwork_10 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_10_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_10_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_10_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_10_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_10_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_10_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_10_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_10_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_10_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_10_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_10_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_10_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_10_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_10_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_10_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_10_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_10_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_10_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_10_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_10_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_10_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_10_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_10_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_10_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_10_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_10_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_10_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_10_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_10_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_10_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_10_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_10_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_10_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_10_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_10_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_10_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_10_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_10_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_10_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_10_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_10_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_10_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_10_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_10_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_10_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_10_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_10_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_10_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_10_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_10_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_10_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_10_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_10_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_10_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_10_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_10_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_10_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_10_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_10_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_10_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_10_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_10_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_10_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_10_io_to_mem_bits)
  );
  PENetwork PENetwork_11 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_11_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_11_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_11_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_11_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_11_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_11_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_11_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_11_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_11_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_11_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_11_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_11_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_11_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_11_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_11_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_11_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_11_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_11_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_11_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_11_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_11_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_11_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_11_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_11_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_11_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_11_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_11_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_11_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_11_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_11_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_11_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_11_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_11_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_11_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_11_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_11_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_11_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_11_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_11_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_11_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_11_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_11_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_11_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_11_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_11_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_11_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_11_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_11_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_11_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_11_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_11_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_11_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_11_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_11_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_11_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_11_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_11_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_11_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_11_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_11_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_11_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_11_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_11_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_11_io_to_mem_bits)
  );
  PENetwork PENetwork_12 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_12_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_12_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_12_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_12_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_12_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_12_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_12_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_12_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_12_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_12_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_12_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_12_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_12_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_12_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_12_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_12_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_12_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_12_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_12_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_12_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_12_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_12_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_12_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_12_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_12_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_12_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_12_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_12_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_12_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_12_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_12_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_12_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_12_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_12_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_12_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_12_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_12_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_12_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_12_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_12_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_12_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_12_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_12_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_12_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_12_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_12_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_12_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_12_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_12_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_12_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_12_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_12_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_12_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_12_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_12_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_12_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_12_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_12_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_12_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_12_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_12_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_12_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_12_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_12_io_to_mem_bits)
  );
  PENetwork PENetwork_13 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_13_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_13_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_13_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_13_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_13_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_13_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_13_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_13_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_13_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_13_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_13_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_13_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_13_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_13_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_13_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_13_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_13_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_13_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_13_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_13_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_13_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_13_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_13_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_13_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_13_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_13_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_13_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_13_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_13_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_13_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_13_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_13_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_13_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_13_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_13_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_13_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_13_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_13_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_13_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_13_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_13_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_13_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_13_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_13_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_13_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_13_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_13_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_13_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_13_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_13_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_13_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_13_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_13_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_13_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_13_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_13_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_13_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_13_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_13_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_13_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_13_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_13_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_13_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_13_io_to_mem_bits)
  );
  PENetwork PENetwork_14 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_14_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_14_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_14_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_14_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_14_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_14_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_14_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_14_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_14_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_14_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_14_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_14_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_14_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_14_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_14_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_14_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_14_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_14_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_14_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_14_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_14_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_14_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_14_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_14_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_14_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_14_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_14_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_14_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_14_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_14_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_14_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_14_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_14_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_14_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_14_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_14_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_14_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_14_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_14_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_14_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_14_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_14_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_14_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_14_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_14_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_14_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_14_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_14_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_14_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_14_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_14_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_14_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_14_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_14_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_14_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_14_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_14_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_14_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_14_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_14_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_14_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_14_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_14_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_14_io_to_mem_bits)
  );
  PENetwork PENetwork_15 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_15_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_15_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_15_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_15_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_15_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_15_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_15_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_15_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_15_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_15_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_15_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_15_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_15_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_15_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_15_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_15_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_15_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_15_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_15_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_15_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_15_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_15_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_15_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_15_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_15_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_15_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_15_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_15_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_15_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_15_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_15_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_15_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_15_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_15_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_15_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_15_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_15_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_15_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_15_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_15_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_15_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_15_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_15_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_15_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_15_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_15_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_15_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_15_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_15_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_15_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_15_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_15_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_15_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_15_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_15_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_15_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_15_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_15_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_15_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_15_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_15_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_15_io_to_pes_15_out_bits),
    .io_to_mem_valid(PENetwork_15_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_15_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_16 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_16_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_16_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_16_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_16_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_16_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_16_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_16_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_16_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_16_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_16_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_16_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_16_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_16_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_16_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_16_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_16_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_16_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_16_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_16_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_16_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_16_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_16_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_16_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_16_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_16_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_16_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_16_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_16_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_16_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_16_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_16_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_16_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_16_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_16_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_16_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_16_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_16_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_16_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_16_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_16_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_16_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_16_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_16_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_16_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_16_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_16_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_16_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_16_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_16_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_16_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_16_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_16_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_16_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_16_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_16_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_16_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_16_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_16_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_16_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_16_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_16_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_16_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_16_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_16_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_17 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_17_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_17_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_17_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_17_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_17_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_17_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_17_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_17_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_17_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_17_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_17_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_17_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_17_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_17_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_17_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_17_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_17_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_17_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_17_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_17_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_17_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_17_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_17_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_17_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_17_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_17_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_17_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_17_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_17_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_17_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_17_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_17_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_17_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_17_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_17_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_17_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_17_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_17_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_17_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_17_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_17_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_17_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_17_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_17_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_17_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_17_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_17_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_17_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_17_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_17_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_17_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_17_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_17_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_17_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_17_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_17_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_17_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_17_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_17_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_17_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_17_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_17_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_17_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_17_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_18 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_18_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_18_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_18_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_18_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_18_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_18_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_18_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_18_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_18_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_18_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_18_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_18_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_18_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_18_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_18_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_18_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_18_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_18_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_18_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_18_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_18_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_18_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_18_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_18_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_18_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_18_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_18_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_18_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_18_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_18_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_18_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_18_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_18_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_18_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_18_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_18_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_18_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_18_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_18_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_18_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_18_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_18_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_18_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_18_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_18_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_18_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_18_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_18_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_18_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_18_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_18_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_18_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_18_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_18_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_18_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_18_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_18_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_18_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_18_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_18_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_18_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_18_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_18_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_18_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_19 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_19_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_19_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_19_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_19_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_19_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_19_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_19_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_19_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_19_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_19_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_19_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_19_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_19_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_19_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_19_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_19_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_19_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_19_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_19_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_19_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_19_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_19_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_19_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_19_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_19_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_19_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_19_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_19_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_19_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_19_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_19_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_19_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_19_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_19_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_19_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_19_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_19_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_19_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_19_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_19_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_19_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_19_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_19_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_19_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_19_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_19_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_19_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_19_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_19_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_19_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_19_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_19_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_19_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_19_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_19_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_19_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_19_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_19_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_19_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_19_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_19_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_19_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_19_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_19_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_20 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_20_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_20_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_20_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_20_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_20_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_20_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_20_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_20_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_20_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_20_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_20_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_20_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_20_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_20_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_20_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_20_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_20_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_20_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_20_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_20_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_20_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_20_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_20_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_20_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_20_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_20_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_20_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_20_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_20_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_20_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_20_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_20_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_20_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_20_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_20_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_20_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_20_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_20_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_20_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_20_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_20_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_20_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_20_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_20_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_20_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_20_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_20_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_20_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_20_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_20_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_20_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_20_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_20_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_20_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_20_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_20_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_20_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_20_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_20_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_20_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_20_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_20_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_20_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_20_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_21 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_21_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_21_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_21_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_21_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_21_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_21_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_21_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_21_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_21_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_21_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_21_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_21_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_21_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_21_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_21_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_21_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_21_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_21_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_21_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_21_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_21_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_21_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_21_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_21_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_21_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_21_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_21_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_21_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_21_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_21_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_21_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_21_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_21_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_21_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_21_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_21_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_21_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_21_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_21_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_21_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_21_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_21_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_21_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_21_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_21_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_21_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_21_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_21_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_21_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_21_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_21_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_21_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_21_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_21_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_21_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_21_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_21_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_21_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_21_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_21_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_21_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_21_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_21_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_21_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_22 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_22_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_22_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_22_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_22_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_22_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_22_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_22_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_22_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_22_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_22_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_22_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_22_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_22_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_22_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_22_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_22_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_22_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_22_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_22_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_22_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_22_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_22_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_22_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_22_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_22_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_22_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_22_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_22_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_22_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_22_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_22_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_22_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_22_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_22_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_22_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_22_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_22_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_22_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_22_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_22_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_22_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_22_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_22_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_22_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_22_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_22_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_22_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_22_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_22_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_22_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_22_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_22_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_22_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_22_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_22_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_22_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_22_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_22_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_22_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_22_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_22_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_22_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_22_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_22_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_23 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_23_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_23_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_23_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_23_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_23_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_23_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_23_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_23_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_23_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_23_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_23_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_23_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_23_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_23_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_23_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_23_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_23_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_23_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_23_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_23_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_23_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_23_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_23_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_23_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_23_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_23_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_23_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_23_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_23_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_23_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_23_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_23_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_23_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_23_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_23_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_23_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_23_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_23_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_23_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_23_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_23_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_23_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_23_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_23_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_23_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_23_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_23_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_23_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_23_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_23_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_23_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_23_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_23_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_23_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_23_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_23_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_23_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_23_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_23_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_23_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_23_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_23_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_23_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_23_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_24 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_24_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_24_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_24_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_24_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_24_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_24_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_24_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_24_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_24_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_24_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_24_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_24_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_24_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_24_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_24_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_24_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_24_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_24_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_24_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_24_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_24_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_24_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_24_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_24_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_24_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_24_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_24_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_24_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_24_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_24_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_24_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_24_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_24_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_24_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_24_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_24_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_24_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_24_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_24_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_24_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_24_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_24_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_24_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_24_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_24_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_24_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_24_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_24_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_24_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_24_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_24_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_24_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_24_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_24_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_24_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_24_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_24_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_24_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_24_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_24_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_24_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_24_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_24_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_24_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_25 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_25_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_25_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_25_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_25_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_25_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_25_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_25_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_25_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_25_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_25_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_25_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_25_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_25_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_25_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_25_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_25_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_25_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_25_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_25_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_25_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_25_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_25_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_25_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_25_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_25_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_25_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_25_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_25_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_25_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_25_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_25_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_25_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_25_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_25_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_25_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_25_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_25_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_25_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_25_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_25_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_25_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_25_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_25_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_25_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_25_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_25_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_25_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_25_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_25_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_25_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_25_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_25_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_25_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_25_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_25_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_25_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_25_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_25_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_25_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_25_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_25_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_25_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_25_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_25_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_26 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_26_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_26_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_26_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_26_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_26_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_26_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_26_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_26_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_26_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_26_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_26_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_26_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_26_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_26_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_26_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_26_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_26_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_26_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_26_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_26_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_26_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_26_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_26_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_26_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_26_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_26_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_26_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_26_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_26_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_26_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_26_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_26_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_26_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_26_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_26_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_26_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_26_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_26_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_26_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_26_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_26_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_26_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_26_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_26_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_26_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_26_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_26_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_26_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_26_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_26_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_26_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_26_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_26_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_26_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_26_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_26_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_26_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_26_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_26_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_26_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_26_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_26_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_26_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_26_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_27 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_27_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_27_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_27_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_27_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_27_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_27_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_27_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_27_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_27_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_27_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_27_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_27_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_27_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_27_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_27_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_27_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_27_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_27_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_27_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_27_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_27_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_27_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_27_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_27_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_27_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_27_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_27_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_27_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_27_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_27_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_27_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_27_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_27_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_27_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_27_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_27_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_27_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_27_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_27_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_27_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_27_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_27_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_27_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_27_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_27_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_27_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_27_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_27_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_27_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_27_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_27_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_27_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_27_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_27_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_27_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_27_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_27_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_27_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_27_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_27_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_27_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_27_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_27_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_27_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_28 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_28_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_28_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_28_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_28_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_28_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_28_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_28_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_28_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_28_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_28_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_28_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_28_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_28_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_28_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_28_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_28_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_28_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_28_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_28_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_28_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_28_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_28_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_28_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_28_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_28_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_28_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_28_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_28_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_28_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_28_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_28_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_28_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_28_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_28_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_28_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_28_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_28_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_28_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_28_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_28_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_28_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_28_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_28_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_28_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_28_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_28_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_28_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_28_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_28_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_28_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_28_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_28_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_28_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_28_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_28_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_28_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_28_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_28_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_28_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_28_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_28_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_28_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_28_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_28_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_29 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_29_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_29_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_29_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_29_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_29_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_29_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_29_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_29_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_29_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_29_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_29_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_29_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_29_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_29_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_29_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_29_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_29_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_29_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_29_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_29_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_29_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_29_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_29_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_29_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_29_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_29_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_29_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_29_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_29_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_29_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_29_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_29_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_29_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_29_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_29_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_29_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_29_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_29_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_29_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_29_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_29_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_29_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_29_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_29_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_29_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_29_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_29_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_29_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_29_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_29_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_29_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_29_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_29_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_29_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_29_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_29_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_29_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_29_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_29_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_29_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_29_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_29_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_29_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_29_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_30 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_30_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_30_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_30_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_30_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_30_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_30_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_30_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_30_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_30_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_30_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_30_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_30_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_30_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_30_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_30_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_30_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_30_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_30_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_30_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_30_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_30_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_30_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_30_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_30_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_30_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_30_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_30_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_30_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_30_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_30_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_30_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_30_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_30_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_30_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_30_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_30_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_30_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_30_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_30_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_30_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_30_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_30_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_30_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_30_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_30_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_30_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_30_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_30_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_30_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_30_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_30_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_30_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_30_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_30_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_30_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_30_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_30_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_30_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_30_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_30_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_30_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_30_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_30_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_30_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_31 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_31_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_31_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_31_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_31_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_31_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_31_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_31_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_31_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_31_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_31_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_31_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_31_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_31_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_31_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_31_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_31_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_31_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_31_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_31_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_31_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_31_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_31_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_31_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_31_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_31_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_31_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_31_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_31_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_31_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_31_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_31_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_31_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_31_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_31_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_31_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_31_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_31_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_31_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_31_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_31_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_31_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_31_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_31_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_31_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_31_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_31_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_31_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_31_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_31_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_31_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_31_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_31_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_31_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_31_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_31_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_31_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_31_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_31_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_31_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_31_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_31_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_31_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_31_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_31_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_32 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_32_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_32_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_32_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_32_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_32_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_32_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_32_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_32_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_32_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_32_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_32_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_32_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_32_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_32_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_32_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_32_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_32_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_32_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_32_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_32_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_32_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_32_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_32_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_32_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_32_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_32_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_32_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_32_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_32_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_32_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_32_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_32_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_32_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_32_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_32_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_32_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_32_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_32_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_32_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_32_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_32_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_32_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_32_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_32_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_32_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_32_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_32_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_32_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_32_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_32_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_32_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_32_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_32_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_32_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_32_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_32_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_32_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_32_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_32_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_32_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_32_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_32_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_32_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_32_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_33 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_33_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_33_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_33_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_33_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_33_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_33_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_33_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_33_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_33_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_33_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_33_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_33_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_33_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_33_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_33_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_33_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_33_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_33_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_33_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_33_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_33_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_33_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_33_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_33_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_33_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_33_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_33_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_33_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_33_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_33_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_33_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_33_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_33_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_33_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_33_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_33_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_33_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_33_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_33_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_33_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_33_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_33_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_33_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_33_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_33_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_33_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_33_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_33_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_33_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_33_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_33_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_33_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_33_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_33_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_33_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_33_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_33_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_33_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_33_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_33_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_33_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_33_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_33_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_33_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_34 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_34_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_34_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_34_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_34_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_34_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_34_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_34_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_34_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_34_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_34_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_34_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_34_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_34_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_34_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_34_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_34_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_34_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_34_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_34_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_34_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_34_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_34_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_34_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_34_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_34_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_34_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_34_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_34_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_34_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_34_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_34_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_34_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_34_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_34_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_34_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_34_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_34_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_34_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_34_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_34_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_34_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_34_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_34_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_34_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_34_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_34_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_34_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_34_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_34_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_34_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_34_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_34_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_34_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_34_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_34_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_34_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_34_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_34_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_34_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_34_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_34_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_34_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_34_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_34_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_35 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_35_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_35_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_35_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_35_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_35_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_35_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_35_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_35_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_35_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_35_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_35_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_35_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_35_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_35_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_35_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_35_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_35_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_35_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_35_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_35_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_35_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_35_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_35_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_35_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_35_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_35_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_35_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_35_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_35_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_35_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_35_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_35_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_35_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_35_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_35_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_35_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_35_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_35_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_35_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_35_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_35_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_35_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_35_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_35_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_35_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_35_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_35_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_35_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_35_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_35_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_35_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_35_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_35_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_35_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_35_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_35_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_35_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_35_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_35_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_35_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_35_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_35_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_35_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_35_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_36 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_36_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_36_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_36_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_36_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_36_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_36_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_36_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_36_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_36_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_36_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_36_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_36_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_36_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_36_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_36_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_36_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_36_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_36_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_36_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_36_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_36_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_36_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_36_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_36_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_36_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_36_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_36_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_36_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_36_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_36_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_36_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_36_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_36_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_36_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_36_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_36_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_36_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_36_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_36_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_36_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_36_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_36_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_36_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_36_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_36_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_36_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_36_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_36_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_36_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_36_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_36_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_36_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_36_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_36_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_36_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_36_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_36_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_36_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_36_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_36_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_36_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_36_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_36_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_36_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_37 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_37_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_37_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_37_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_37_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_37_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_37_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_37_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_37_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_37_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_37_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_37_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_37_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_37_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_37_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_37_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_37_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_37_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_37_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_37_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_37_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_37_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_37_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_37_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_37_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_37_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_37_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_37_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_37_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_37_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_37_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_37_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_37_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_37_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_37_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_37_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_37_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_37_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_37_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_37_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_37_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_37_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_37_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_37_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_37_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_37_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_37_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_37_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_37_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_37_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_37_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_37_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_37_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_37_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_37_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_37_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_37_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_37_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_37_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_37_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_37_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_37_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_37_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_37_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_37_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_38 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_38_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_38_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_38_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_38_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_38_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_38_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_38_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_38_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_38_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_38_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_38_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_38_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_38_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_38_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_38_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_38_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_38_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_38_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_38_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_38_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_38_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_38_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_38_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_38_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_38_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_38_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_38_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_38_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_38_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_38_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_38_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_38_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_38_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_38_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_38_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_38_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_38_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_38_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_38_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_38_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_38_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_38_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_38_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_38_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_38_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_38_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_38_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_38_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_38_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_38_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_38_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_38_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_38_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_38_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_38_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_38_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_38_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_38_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_38_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_38_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_38_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_38_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_38_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_38_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_39 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_39_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_39_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_39_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_39_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_39_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_39_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_39_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_39_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_39_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_39_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_39_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_39_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_39_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_39_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_39_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_39_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_39_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_39_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_39_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_39_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_39_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_39_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_39_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_39_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_39_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_39_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_39_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_39_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_39_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_39_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_39_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_39_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_39_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_39_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_39_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_39_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_39_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_39_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_39_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_39_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_39_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_39_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_39_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_39_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_39_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_39_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_39_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_39_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_39_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_39_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_39_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_39_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_39_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_39_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_39_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_39_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_39_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_39_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_39_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_39_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_39_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_39_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_39_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_39_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_40 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_40_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_40_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_40_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_40_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_40_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_40_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_40_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_40_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_40_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_40_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_40_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_40_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_40_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_40_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_40_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_40_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_40_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_40_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_40_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_40_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_40_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_40_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_40_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_40_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_40_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_40_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_40_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_40_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_40_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_40_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_40_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_40_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_40_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_40_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_40_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_40_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_40_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_40_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_40_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_40_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_40_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_40_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_40_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_40_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_40_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_40_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_40_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_40_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_40_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_40_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_40_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_40_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_40_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_40_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_40_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_40_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_40_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_40_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_40_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_40_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_40_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_40_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_40_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_40_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_41 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_41_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_41_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_41_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_41_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_41_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_41_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_41_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_41_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_41_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_41_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_41_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_41_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_41_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_41_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_41_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_41_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_41_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_41_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_41_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_41_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_41_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_41_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_41_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_41_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_41_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_41_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_41_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_41_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_41_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_41_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_41_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_41_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_41_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_41_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_41_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_41_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_41_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_41_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_41_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_41_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_41_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_41_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_41_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_41_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_41_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_41_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_41_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_41_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_41_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_41_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_41_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_41_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_41_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_41_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_41_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_41_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_41_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_41_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_41_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_41_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_41_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_41_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_41_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_41_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_42 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_42_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_42_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_42_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_42_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_42_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_42_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_42_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_42_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_42_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_42_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_42_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_42_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_42_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_42_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_42_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_42_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_42_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_42_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_42_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_42_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_42_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_42_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_42_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_42_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_42_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_42_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_42_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_42_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_42_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_42_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_42_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_42_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_42_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_42_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_42_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_42_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_42_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_42_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_42_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_42_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_42_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_42_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_42_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_42_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_42_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_42_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_42_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_42_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_42_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_42_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_42_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_42_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_42_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_42_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_42_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_42_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_42_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_42_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_42_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_42_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_42_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_42_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_42_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_42_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_43 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_43_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_43_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_43_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_43_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_43_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_43_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_43_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_43_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_43_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_43_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_43_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_43_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_43_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_43_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_43_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_43_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_43_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_43_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_43_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_43_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_43_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_43_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_43_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_43_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_43_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_43_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_43_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_43_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_43_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_43_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_43_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_43_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_43_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_43_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_43_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_43_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_43_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_43_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_43_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_43_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_43_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_43_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_43_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_43_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_43_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_43_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_43_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_43_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_43_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_43_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_43_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_43_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_43_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_43_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_43_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_43_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_43_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_43_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_43_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_43_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_43_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_43_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_43_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_43_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_44 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_44_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_44_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_44_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_44_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_44_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_44_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_44_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_44_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_44_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_44_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_44_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_44_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_44_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_44_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_44_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_44_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_44_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_44_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_44_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_44_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_44_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_44_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_44_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_44_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_44_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_44_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_44_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_44_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_44_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_44_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_44_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_44_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_44_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_44_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_44_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_44_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_44_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_44_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_44_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_44_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_44_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_44_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_44_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_44_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_44_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_44_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_44_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_44_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_44_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_44_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_44_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_44_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_44_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_44_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_44_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_44_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_44_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_44_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_44_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_44_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_44_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_44_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_44_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_44_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_45 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_45_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_45_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_45_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_45_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_45_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_45_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_45_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_45_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_45_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_45_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_45_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_45_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_45_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_45_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_45_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_45_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_45_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_45_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_45_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_45_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_45_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_45_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_45_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_45_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_45_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_45_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_45_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_45_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_45_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_45_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_45_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_45_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_45_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_45_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_45_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_45_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_45_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_45_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_45_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_45_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_45_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_45_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_45_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_45_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_45_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_45_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_45_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_45_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_45_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_45_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_45_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_45_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_45_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_45_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_45_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_45_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_45_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_45_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_45_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_45_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_45_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_45_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_45_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_45_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_46 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_46_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_46_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_46_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_46_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_46_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_46_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_46_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_46_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_46_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_46_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_46_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_46_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_46_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_46_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_46_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_46_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_46_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_46_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_46_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_46_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_46_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_46_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_46_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_46_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_46_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_46_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_46_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_46_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_46_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_46_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_46_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_46_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_46_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_46_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_46_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_46_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_46_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_46_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_46_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_46_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_46_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_46_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_46_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_46_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_46_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_46_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_46_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_46_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_46_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_46_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_46_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_46_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_46_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_46_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_46_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_46_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_46_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_46_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_46_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_46_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_46_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_46_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_46_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_46_io_to_mem_bits)
  );
  PENetwork_16 PENetwork_47 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_47_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_47_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_47_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_47_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_47_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_47_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_47_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_47_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_47_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_47_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_47_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_47_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_47_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_47_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_47_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_47_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_47_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_47_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_47_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_47_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_47_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_47_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_47_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_47_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_47_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_47_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_47_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_47_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_47_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_47_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_47_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_47_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_47_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_47_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_47_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_47_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_47_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_47_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_47_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_47_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_47_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_47_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_47_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_47_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_47_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_47_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_47_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_47_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_47_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_47_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_47_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_47_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_47_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_47_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_47_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_47_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_47_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_47_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_47_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_47_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_47_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_47_io_to_pes_15_in_bits),
    .io_to_mem_valid(PENetwork_47_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_47_io_to_mem_bits)
  );
  MemController MemController ( // @[pearray.scala 212:15]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_rd_valid(MemController_io_rd_valid),
    .io_wr_valid(MemController_io_wr_valid),
    .io_rd_data_valid(MemController_io_rd_data_valid),
    .io_rd_data_bits(MemController_io_rd_data_bits),
    .io_wr_data_valid(MemController_io_wr_data_valid),
    .io_wr_data_bits(MemController_io_wr_data_bits)
  );
  MemController MemController_1 ( // @[pearray.scala 212:15]
    .clock(MemController_1_clock),
    .reset(MemController_1_reset),
    .io_rd_valid(MemController_1_io_rd_valid),
    .io_wr_valid(MemController_1_io_wr_valid),
    .io_rd_data_valid(MemController_1_io_rd_data_valid),
    .io_rd_data_bits(MemController_1_io_rd_data_bits),
    .io_wr_data_valid(MemController_1_io_wr_data_valid),
    .io_wr_data_bits(MemController_1_io_wr_data_bits)
  );
  MemController MemController_2 ( // @[pearray.scala 212:15]
    .clock(MemController_2_clock),
    .reset(MemController_2_reset),
    .io_rd_valid(MemController_2_io_rd_valid),
    .io_wr_valid(MemController_2_io_wr_valid),
    .io_rd_data_valid(MemController_2_io_rd_data_valid),
    .io_rd_data_bits(MemController_2_io_rd_data_bits),
    .io_wr_data_valid(MemController_2_io_wr_data_valid),
    .io_wr_data_bits(MemController_2_io_wr_data_bits)
  );
  MemController MemController_3 ( // @[pearray.scala 212:15]
    .clock(MemController_3_clock),
    .reset(MemController_3_reset),
    .io_rd_valid(MemController_3_io_rd_valid),
    .io_wr_valid(MemController_3_io_wr_valid),
    .io_rd_data_valid(MemController_3_io_rd_data_valid),
    .io_rd_data_bits(MemController_3_io_rd_data_bits),
    .io_wr_data_valid(MemController_3_io_wr_data_valid),
    .io_wr_data_bits(MemController_3_io_wr_data_bits)
  );
  MemController MemController_4 ( // @[pearray.scala 212:15]
    .clock(MemController_4_clock),
    .reset(MemController_4_reset),
    .io_rd_valid(MemController_4_io_rd_valid),
    .io_wr_valid(MemController_4_io_wr_valid),
    .io_rd_data_valid(MemController_4_io_rd_data_valid),
    .io_rd_data_bits(MemController_4_io_rd_data_bits),
    .io_wr_data_valid(MemController_4_io_wr_data_valid),
    .io_wr_data_bits(MemController_4_io_wr_data_bits)
  );
  MemController MemController_5 ( // @[pearray.scala 212:15]
    .clock(MemController_5_clock),
    .reset(MemController_5_reset),
    .io_rd_valid(MemController_5_io_rd_valid),
    .io_wr_valid(MemController_5_io_wr_valid),
    .io_rd_data_valid(MemController_5_io_rd_data_valid),
    .io_rd_data_bits(MemController_5_io_rd_data_bits),
    .io_wr_data_valid(MemController_5_io_wr_data_valid),
    .io_wr_data_bits(MemController_5_io_wr_data_bits)
  );
  MemController MemController_6 ( // @[pearray.scala 212:15]
    .clock(MemController_6_clock),
    .reset(MemController_6_reset),
    .io_rd_valid(MemController_6_io_rd_valid),
    .io_wr_valid(MemController_6_io_wr_valid),
    .io_rd_data_valid(MemController_6_io_rd_data_valid),
    .io_rd_data_bits(MemController_6_io_rd_data_bits),
    .io_wr_data_valid(MemController_6_io_wr_data_valid),
    .io_wr_data_bits(MemController_6_io_wr_data_bits)
  );
  MemController MemController_7 ( // @[pearray.scala 212:15]
    .clock(MemController_7_clock),
    .reset(MemController_7_reset),
    .io_rd_valid(MemController_7_io_rd_valid),
    .io_wr_valid(MemController_7_io_wr_valid),
    .io_rd_data_valid(MemController_7_io_rd_data_valid),
    .io_rd_data_bits(MemController_7_io_rd_data_bits),
    .io_wr_data_valid(MemController_7_io_wr_data_valid),
    .io_wr_data_bits(MemController_7_io_wr_data_bits)
  );
  MemController MemController_8 ( // @[pearray.scala 212:15]
    .clock(MemController_8_clock),
    .reset(MemController_8_reset),
    .io_rd_valid(MemController_8_io_rd_valid),
    .io_wr_valid(MemController_8_io_wr_valid),
    .io_rd_data_valid(MemController_8_io_rd_data_valid),
    .io_rd_data_bits(MemController_8_io_rd_data_bits),
    .io_wr_data_valid(MemController_8_io_wr_data_valid),
    .io_wr_data_bits(MemController_8_io_wr_data_bits)
  );
  MemController MemController_9 ( // @[pearray.scala 212:15]
    .clock(MemController_9_clock),
    .reset(MemController_9_reset),
    .io_rd_valid(MemController_9_io_rd_valid),
    .io_wr_valid(MemController_9_io_wr_valid),
    .io_rd_data_valid(MemController_9_io_rd_data_valid),
    .io_rd_data_bits(MemController_9_io_rd_data_bits),
    .io_wr_data_valid(MemController_9_io_wr_data_valid),
    .io_wr_data_bits(MemController_9_io_wr_data_bits)
  );
  MemController MemController_10 ( // @[pearray.scala 212:15]
    .clock(MemController_10_clock),
    .reset(MemController_10_reset),
    .io_rd_valid(MemController_10_io_rd_valid),
    .io_wr_valid(MemController_10_io_wr_valid),
    .io_rd_data_valid(MemController_10_io_rd_data_valid),
    .io_rd_data_bits(MemController_10_io_rd_data_bits),
    .io_wr_data_valid(MemController_10_io_wr_data_valid),
    .io_wr_data_bits(MemController_10_io_wr_data_bits)
  );
  MemController MemController_11 ( // @[pearray.scala 212:15]
    .clock(MemController_11_clock),
    .reset(MemController_11_reset),
    .io_rd_valid(MemController_11_io_rd_valid),
    .io_wr_valid(MemController_11_io_wr_valid),
    .io_rd_data_valid(MemController_11_io_rd_data_valid),
    .io_rd_data_bits(MemController_11_io_rd_data_bits),
    .io_wr_data_valid(MemController_11_io_wr_data_valid),
    .io_wr_data_bits(MemController_11_io_wr_data_bits)
  );
  MemController MemController_12 ( // @[pearray.scala 212:15]
    .clock(MemController_12_clock),
    .reset(MemController_12_reset),
    .io_rd_valid(MemController_12_io_rd_valid),
    .io_wr_valid(MemController_12_io_wr_valid),
    .io_rd_data_valid(MemController_12_io_rd_data_valid),
    .io_rd_data_bits(MemController_12_io_rd_data_bits),
    .io_wr_data_valid(MemController_12_io_wr_data_valid),
    .io_wr_data_bits(MemController_12_io_wr_data_bits)
  );
  MemController MemController_13 ( // @[pearray.scala 212:15]
    .clock(MemController_13_clock),
    .reset(MemController_13_reset),
    .io_rd_valid(MemController_13_io_rd_valid),
    .io_wr_valid(MemController_13_io_wr_valid),
    .io_rd_data_valid(MemController_13_io_rd_data_valid),
    .io_rd_data_bits(MemController_13_io_rd_data_bits),
    .io_wr_data_valid(MemController_13_io_wr_data_valid),
    .io_wr_data_bits(MemController_13_io_wr_data_bits)
  );
  MemController MemController_14 ( // @[pearray.scala 212:15]
    .clock(MemController_14_clock),
    .reset(MemController_14_reset),
    .io_rd_valid(MemController_14_io_rd_valid),
    .io_wr_valid(MemController_14_io_wr_valid),
    .io_rd_data_valid(MemController_14_io_rd_data_valid),
    .io_rd_data_bits(MemController_14_io_rd_data_bits),
    .io_wr_data_valid(MemController_14_io_wr_data_valid),
    .io_wr_data_bits(MemController_14_io_wr_data_bits)
  );
  MemController MemController_15 ( // @[pearray.scala 212:15]
    .clock(MemController_15_clock),
    .reset(MemController_15_reset),
    .io_rd_valid(MemController_15_io_rd_valid),
    .io_wr_valid(MemController_15_io_wr_valid),
    .io_rd_data_valid(MemController_15_io_rd_data_valid),
    .io_rd_data_bits(MemController_15_io_rd_data_bits),
    .io_wr_data_valid(MemController_15_io_wr_data_valid),
    .io_wr_data_bits(MemController_15_io_wr_data_bits)
  );
  MemController_16 MemController_16 ( // @[pearray.scala 210:15]
    .clock(MemController_16_clock),
    .reset(MemController_16_reset),
    .io_rd_valid(MemController_16_io_rd_valid),
    .io_wr_valid(MemController_16_io_wr_valid),
    .io_rd_data_valid(MemController_16_io_rd_data_valid),
    .io_rd_data_bits(MemController_16_io_rd_data_bits),
    .io_wr_data_valid(MemController_16_io_wr_data_valid),
    .io_wr_data_bits(MemController_16_io_wr_data_bits)
  );
  MemController_16 MemController_17 ( // @[pearray.scala 210:15]
    .clock(MemController_17_clock),
    .reset(MemController_17_reset),
    .io_rd_valid(MemController_17_io_rd_valid),
    .io_wr_valid(MemController_17_io_wr_valid),
    .io_rd_data_valid(MemController_17_io_rd_data_valid),
    .io_rd_data_bits(MemController_17_io_rd_data_bits),
    .io_wr_data_valid(MemController_17_io_wr_data_valid),
    .io_wr_data_bits(MemController_17_io_wr_data_bits)
  );
  MemController_16 MemController_18 ( // @[pearray.scala 210:15]
    .clock(MemController_18_clock),
    .reset(MemController_18_reset),
    .io_rd_valid(MemController_18_io_rd_valid),
    .io_wr_valid(MemController_18_io_wr_valid),
    .io_rd_data_valid(MemController_18_io_rd_data_valid),
    .io_rd_data_bits(MemController_18_io_rd_data_bits),
    .io_wr_data_valid(MemController_18_io_wr_data_valid),
    .io_wr_data_bits(MemController_18_io_wr_data_bits)
  );
  MemController_16 MemController_19 ( // @[pearray.scala 210:15]
    .clock(MemController_19_clock),
    .reset(MemController_19_reset),
    .io_rd_valid(MemController_19_io_rd_valid),
    .io_wr_valid(MemController_19_io_wr_valid),
    .io_rd_data_valid(MemController_19_io_rd_data_valid),
    .io_rd_data_bits(MemController_19_io_rd_data_bits),
    .io_wr_data_valid(MemController_19_io_wr_data_valid),
    .io_wr_data_bits(MemController_19_io_wr_data_bits)
  );
  MemController_16 MemController_20 ( // @[pearray.scala 210:15]
    .clock(MemController_20_clock),
    .reset(MemController_20_reset),
    .io_rd_valid(MemController_20_io_rd_valid),
    .io_wr_valid(MemController_20_io_wr_valid),
    .io_rd_data_valid(MemController_20_io_rd_data_valid),
    .io_rd_data_bits(MemController_20_io_rd_data_bits),
    .io_wr_data_valid(MemController_20_io_wr_data_valid),
    .io_wr_data_bits(MemController_20_io_wr_data_bits)
  );
  MemController_16 MemController_21 ( // @[pearray.scala 210:15]
    .clock(MemController_21_clock),
    .reset(MemController_21_reset),
    .io_rd_valid(MemController_21_io_rd_valid),
    .io_wr_valid(MemController_21_io_wr_valid),
    .io_rd_data_valid(MemController_21_io_rd_data_valid),
    .io_rd_data_bits(MemController_21_io_rd_data_bits),
    .io_wr_data_valid(MemController_21_io_wr_data_valid),
    .io_wr_data_bits(MemController_21_io_wr_data_bits)
  );
  MemController_16 MemController_22 ( // @[pearray.scala 210:15]
    .clock(MemController_22_clock),
    .reset(MemController_22_reset),
    .io_rd_valid(MemController_22_io_rd_valid),
    .io_wr_valid(MemController_22_io_wr_valid),
    .io_rd_data_valid(MemController_22_io_rd_data_valid),
    .io_rd_data_bits(MemController_22_io_rd_data_bits),
    .io_wr_data_valid(MemController_22_io_wr_data_valid),
    .io_wr_data_bits(MemController_22_io_wr_data_bits)
  );
  MemController_16 MemController_23 ( // @[pearray.scala 210:15]
    .clock(MemController_23_clock),
    .reset(MemController_23_reset),
    .io_rd_valid(MemController_23_io_rd_valid),
    .io_wr_valid(MemController_23_io_wr_valid),
    .io_rd_data_valid(MemController_23_io_rd_data_valid),
    .io_rd_data_bits(MemController_23_io_rd_data_bits),
    .io_wr_data_valid(MemController_23_io_wr_data_valid),
    .io_wr_data_bits(MemController_23_io_wr_data_bits)
  );
  MemController_16 MemController_24 ( // @[pearray.scala 210:15]
    .clock(MemController_24_clock),
    .reset(MemController_24_reset),
    .io_rd_valid(MemController_24_io_rd_valid),
    .io_wr_valid(MemController_24_io_wr_valid),
    .io_rd_data_valid(MemController_24_io_rd_data_valid),
    .io_rd_data_bits(MemController_24_io_rd_data_bits),
    .io_wr_data_valid(MemController_24_io_wr_data_valid),
    .io_wr_data_bits(MemController_24_io_wr_data_bits)
  );
  MemController_16 MemController_25 ( // @[pearray.scala 210:15]
    .clock(MemController_25_clock),
    .reset(MemController_25_reset),
    .io_rd_valid(MemController_25_io_rd_valid),
    .io_wr_valid(MemController_25_io_wr_valid),
    .io_rd_data_valid(MemController_25_io_rd_data_valid),
    .io_rd_data_bits(MemController_25_io_rd_data_bits),
    .io_wr_data_valid(MemController_25_io_wr_data_valid),
    .io_wr_data_bits(MemController_25_io_wr_data_bits)
  );
  MemController_16 MemController_26 ( // @[pearray.scala 210:15]
    .clock(MemController_26_clock),
    .reset(MemController_26_reset),
    .io_rd_valid(MemController_26_io_rd_valid),
    .io_wr_valid(MemController_26_io_wr_valid),
    .io_rd_data_valid(MemController_26_io_rd_data_valid),
    .io_rd_data_bits(MemController_26_io_rd_data_bits),
    .io_wr_data_valid(MemController_26_io_wr_data_valid),
    .io_wr_data_bits(MemController_26_io_wr_data_bits)
  );
  MemController_16 MemController_27 ( // @[pearray.scala 210:15]
    .clock(MemController_27_clock),
    .reset(MemController_27_reset),
    .io_rd_valid(MemController_27_io_rd_valid),
    .io_wr_valid(MemController_27_io_wr_valid),
    .io_rd_data_valid(MemController_27_io_rd_data_valid),
    .io_rd_data_bits(MemController_27_io_rd_data_bits),
    .io_wr_data_valid(MemController_27_io_wr_data_valid),
    .io_wr_data_bits(MemController_27_io_wr_data_bits)
  );
  MemController_16 MemController_28 ( // @[pearray.scala 210:15]
    .clock(MemController_28_clock),
    .reset(MemController_28_reset),
    .io_rd_valid(MemController_28_io_rd_valid),
    .io_wr_valid(MemController_28_io_wr_valid),
    .io_rd_data_valid(MemController_28_io_rd_data_valid),
    .io_rd_data_bits(MemController_28_io_rd_data_bits),
    .io_wr_data_valid(MemController_28_io_wr_data_valid),
    .io_wr_data_bits(MemController_28_io_wr_data_bits)
  );
  MemController_16 MemController_29 ( // @[pearray.scala 210:15]
    .clock(MemController_29_clock),
    .reset(MemController_29_reset),
    .io_rd_valid(MemController_29_io_rd_valid),
    .io_wr_valid(MemController_29_io_wr_valid),
    .io_rd_data_valid(MemController_29_io_rd_data_valid),
    .io_rd_data_bits(MemController_29_io_rd_data_bits),
    .io_wr_data_valid(MemController_29_io_wr_data_valid),
    .io_wr_data_bits(MemController_29_io_wr_data_bits)
  );
  MemController_16 MemController_30 ( // @[pearray.scala 210:15]
    .clock(MemController_30_clock),
    .reset(MemController_30_reset),
    .io_rd_valid(MemController_30_io_rd_valid),
    .io_wr_valid(MemController_30_io_wr_valid),
    .io_rd_data_valid(MemController_30_io_rd_data_valid),
    .io_rd_data_bits(MemController_30_io_rd_data_bits),
    .io_wr_data_valid(MemController_30_io_wr_data_valid),
    .io_wr_data_bits(MemController_30_io_wr_data_bits)
  );
  MemController_16 MemController_31 ( // @[pearray.scala 210:15]
    .clock(MemController_31_clock),
    .reset(MemController_31_reset),
    .io_rd_valid(MemController_31_io_rd_valid),
    .io_wr_valid(MemController_31_io_wr_valid),
    .io_rd_data_valid(MemController_31_io_rd_data_valid),
    .io_rd_data_bits(MemController_31_io_rd_data_bits),
    .io_wr_data_valid(MemController_31_io_wr_data_valid),
    .io_wr_data_bits(MemController_31_io_wr_data_bits)
  );
  MemController_32 MemController_32 ( // @[pearray.scala 210:15]
    .clock(MemController_32_clock),
    .reset(MemController_32_reset),
    .io_rd_valid(MemController_32_io_rd_valid),
    .io_wr_valid(MemController_32_io_wr_valid),
    .io_rd_data_valid(MemController_32_io_rd_data_valid),
    .io_rd_data_bits(MemController_32_io_rd_data_bits),
    .io_wr_data_valid(MemController_32_io_wr_data_valid),
    .io_wr_data_bits(MemController_32_io_wr_data_bits)
  );
  MemController_32 MemController_33 ( // @[pearray.scala 210:15]
    .clock(MemController_33_clock),
    .reset(MemController_33_reset),
    .io_rd_valid(MemController_33_io_rd_valid),
    .io_wr_valid(MemController_33_io_wr_valid),
    .io_rd_data_valid(MemController_33_io_rd_data_valid),
    .io_rd_data_bits(MemController_33_io_rd_data_bits),
    .io_wr_data_valid(MemController_33_io_wr_data_valid),
    .io_wr_data_bits(MemController_33_io_wr_data_bits)
  );
  MemController_32 MemController_34 ( // @[pearray.scala 210:15]
    .clock(MemController_34_clock),
    .reset(MemController_34_reset),
    .io_rd_valid(MemController_34_io_rd_valid),
    .io_wr_valid(MemController_34_io_wr_valid),
    .io_rd_data_valid(MemController_34_io_rd_data_valid),
    .io_rd_data_bits(MemController_34_io_rd_data_bits),
    .io_wr_data_valid(MemController_34_io_wr_data_valid),
    .io_wr_data_bits(MemController_34_io_wr_data_bits)
  );
  MemController_32 MemController_35 ( // @[pearray.scala 210:15]
    .clock(MemController_35_clock),
    .reset(MemController_35_reset),
    .io_rd_valid(MemController_35_io_rd_valid),
    .io_wr_valid(MemController_35_io_wr_valid),
    .io_rd_data_valid(MemController_35_io_rd_data_valid),
    .io_rd_data_bits(MemController_35_io_rd_data_bits),
    .io_wr_data_valid(MemController_35_io_wr_data_valid),
    .io_wr_data_bits(MemController_35_io_wr_data_bits)
  );
  MemController_32 MemController_36 ( // @[pearray.scala 210:15]
    .clock(MemController_36_clock),
    .reset(MemController_36_reset),
    .io_rd_valid(MemController_36_io_rd_valid),
    .io_wr_valid(MemController_36_io_wr_valid),
    .io_rd_data_valid(MemController_36_io_rd_data_valid),
    .io_rd_data_bits(MemController_36_io_rd_data_bits),
    .io_wr_data_valid(MemController_36_io_wr_data_valid),
    .io_wr_data_bits(MemController_36_io_wr_data_bits)
  );
  MemController_32 MemController_37 ( // @[pearray.scala 210:15]
    .clock(MemController_37_clock),
    .reset(MemController_37_reset),
    .io_rd_valid(MemController_37_io_rd_valid),
    .io_wr_valid(MemController_37_io_wr_valid),
    .io_rd_data_valid(MemController_37_io_rd_data_valid),
    .io_rd_data_bits(MemController_37_io_rd_data_bits),
    .io_wr_data_valid(MemController_37_io_wr_data_valid),
    .io_wr_data_bits(MemController_37_io_wr_data_bits)
  );
  MemController_32 MemController_38 ( // @[pearray.scala 210:15]
    .clock(MemController_38_clock),
    .reset(MemController_38_reset),
    .io_rd_valid(MemController_38_io_rd_valid),
    .io_wr_valid(MemController_38_io_wr_valid),
    .io_rd_data_valid(MemController_38_io_rd_data_valid),
    .io_rd_data_bits(MemController_38_io_rd_data_bits),
    .io_wr_data_valid(MemController_38_io_wr_data_valid),
    .io_wr_data_bits(MemController_38_io_wr_data_bits)
  );
  MemController_32 MemController_39 ( // @[pearray.scala 210:15]
    .clock(MemController_39_clock),
    .reset(MemController_39_reset),
    .io_rd_valid(MemController_39_io_rd_valid),
    .io_wr_valid(MemController_39_io_wr_valid),
    .io_rd_data_valid(MemController_39_io_rd_data_valid),
    .io_rd_data_bits(MemController_39_io_rd_data_bits),
    .io_wr_data_valid(MemController_39_io_wr_data_valid),
    .io_wr_data_bits(MemController_39_io_wr_data_bits)
  );
  MemController_32 MemController_40 ( // @[pearray.scala 210:15]
    .clock(MemController_40_clock),
    .reset(MemController_40_reset),
    .io_rd_valid(MemController_40_io_rd_valid),
    .io_wr_valid(MemController_40_io_wr_valid),
    .io_rd_data_valid(MemController_40_io_rd_data_valid),
    .io_rd_data_bits(MemController_40_io_rd_data_bits),
    .io_wr_data_valid(MemController_40_io_wr_data_valid),
    .io_wr_data_bits(MemController_40_io_wr_data_bits)
  );
  MemController_32 MemController_41 ( // @[pearray.scala 210:15]
    .clock(MemController_41_clock),
    .reset(MemController_41_reset),
    .io_rd_valid(MemController_41_io_rd_valid),
    .io_wr_valid(MemController_41_io_wr_valid),
    .io_rd_data_valid(MemController_41_io_rd_data_valid),
    .io_rd_data_bits(MemController_41_io_rd_data_bits),
    .io_wr_data_valid(MemController_41_io_wr_data_valid),
    .io_wr_data_bits(MemController_41_io_wr_data_bits)
  );
  MemController_32 MemController_42 ( // @[pearray.scala 210:15]
    .clock(MemController_42_clock),
    .reset(MemController_42_reset),
    .io_rd_valid(MemController_42_io_rd_valid),
    .io_wr_valid(MemController_42_io_wr_valid),
    .io_rd_data_valid(MemController_42_io_rd_data_valid),
    .io_rd_data_bits(MemController_42_io_rd_data_bits),
    .io_wr_data_valid(MemController_42_io_wr_data_valid),
    .io_wr_data_bits(MemController_42_io_wr_data_bits)
  );
  MemController_32 MemController_43 ( // @[pearray.scala 210:15]
    .clock(MemController_43_clock),
    .reset(MemController_43_reset),
    .io_rd_valid(MemController_43_io_rd_valid),
    .io_wr_valid(MemController_43_io_wr_valid),
    .io_rd_data_valid(MemController_43_io_rd_data_valid),
    .io_rd_data_bits(MemController_43_io_rd_data_bits),
    .io_wr_data_valid(MemController_43_io_wr_data_valid),
    .io_wr_data_bits(MemController_43_io_wr_data_bits)
  );
  MemController_32 MemController_44 ( // @[pearray.scala 210:15]
    .clock(MemController_44_clock),
    .reset(MemController_44_reset),
    .io_rd_valid(MemController_44_io_rd_valid),
    .io_wr_valid(MemController_44_io_wr_valid),
    .io_rd_data_valid(MemController_44_io_rd_data_valid),
    .io_rd_data_bits(MemController_44_io_rd_data_bits),
    .io_wr_data_valid(MemController_44_io_wr_data_valid),
    .io_wr_data_bits(MemController_44_io_wr_data_bits)
  );
  MemController_32 MemController_45 ( // @[pearray.scala 210:15]
    .clock(MemController_45_clock),
    .reset(MemController_45_reset),
    .io_rd_valid(MemController_45_io_rd_valid),
    .io_wr_valid(MemController_45_io_wr_valid),
    .io_rd_data_valid(MemController_45_io_rd_data_valid),
    .io_rd_data_bits(MemController_45_io_rd_data_bits),
    .io_wr_data_valid(MemController_45_io_wr_data_valid),
    .io_wr_data_bits(MemController_45_io_wr_data_bits)
  );
  MemController_32 MemController_46 ( // @[pearray.scala 210:15]
    .clock(MemController_46_clock),
    .reset(MemController_46_reset),
    .io_rd_valid(MemController_46_io_rd_valid),
    .io_wr_valid(MemController_46_io_wr_valid),
    .io_rd_data_valid(MemController_46_io_rd_data_valid),
    .io_rd_data_bits(MemController_46_io_rd_data_bits),
    .io_wr_data_valid(MemController_46_io_wr_data_valid),
    .io_wr_data_bits(MemController_46_io_wr_data_bits)
  );
  MemController_32 MemController_47 ( // @[pearray.scala 210:15]
    .clock(MemController_47_clock),
    .reset(MemController_47_reset),
    .io_rd_valid(MemController_47_io_rd_valid),
    .io_wr_valid(MemController_47_io_wr_valid),
    .io_rd_data_valid(MemController_47_io_rd_data_valid),
    .io_rd_data_bits(MemController_47_io_rd_data_bits),
    .io_wr_data_valid(MemController_47_io_wr_data_valid),
    .io_wr_data_bits(MemController_47_io_wr_data_bits)
  );
  assign io_data_0_out_0_valid = MemController_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_0_bits = MemController_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_1_valid = MemController_1_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_1_bits = MemController_1_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_2_valid = MemController_2_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_2_bits = MemController_2_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_3_valid = MemController_3_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_3_bits = MemController_3_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_4_valid = MemController_4_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_4_bits = MemController_4_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_5_valid = MemController_5_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_5_bits = MemController_5_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_6_valid = MemController_6_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_6_bits = MemController_6_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_7_valid = MemController_7_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_7_bits = MemController_7_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_8_valid = MemController_8_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_8_bits = MemController_8_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_9_valid = MemController_9_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_9_bits = MemController_9_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_10_valid = MemController_10_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_10_bits = MemController_10_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_11_valid = MemController_11_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_11_bits = MemController_11_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_12_valid = MemController_12_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_12_bits = MemController_12_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_13_valid = MemController_13_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_13_bits = MemController_13_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_14_valid = MemController_14_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_14_bits = MemController_14_io_rd_data_bits; // @[pearray.scala 261:31]
  assign io_data_0_out_15_valid = MemController_15_io_rd_data_valid; // @[pearray.scala 261:31]
  assign io_data_0_out_15_bits = MemController_15_io_rd_data_bits; // @[pearray.scala 261:31]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_exec_valid; // @[pearray.scala 149:16]
  assign PE_clock = clock;
  assign PE_reset = reset;
  assign PE_io_data_2_in_valid = PENetwork_32_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_io_data_2_in_bits = PENetwork_32_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_io_data_1_in_valid = PENetwork_16_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_io_data_1_in_bits = PENetwork_16_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_io_sig_stat2trans = _T_12_3; // @[pearray.scala 184:38]
  assign PE_1_clock = clock;
  assign PE_1_reset = reset;
  assign PE_1_io_data_2_in_valid = PENetwork_33_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_1_io_data_2_in_bits = PENetwork_33_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_1_io_data_1_in_valid = PENetwork_16_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_1_io_data_1_in_bits = PENetwork_16_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_1_io_data_0_in_valid = PENetwork_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_1_io_data_0_in_bits = PENetwork_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_1_io_sig_stat2trans = _T_22_3; // @[pearray.scala 184:38]
  assign PE_2_clock = clock;
  assign PE_2_reset = reset;
  assign PE_2_io_data_2_in_valid = PENetwork_34_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_2_io_data_2_in_bits = PENetwork_34_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_2_io_data_1_in_valid = PENetwork_16_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_2_io_data_1_in_bits = PENetwork_16_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_2_io_data_0_in_valid = PENetwork_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_2_io_data_0_in_bits = PENetwork_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_2_io_sig_stat2trans = _T_32_3; // @[pearray.scala 184:38]
  assign PE_3_clock = clock;
  assign PE_3_reset = reset;
  assign PE_3_io_data_2_in_valid = PENetwork_35_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_3_io_data_2_in_bits = PENetwork_35_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_3_io_data_1_in_valid = PENetwork_16_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_3_io_data_1_in_bits = PENetwork_16_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_3_io_data_0_in_valid = PENetwork_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_3_io_data_0_in_bits = PENetwork_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_3_io_sig_stat2trans = _T_42_3; // @[pearray.scala 184:38]
  assign PE_4_clock = clock;
  assign PE_4_reset = reset;
  assign PE_4_io_data_2_in_valid = PENetwork_36_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_4_io_data_2_in_bits = PENetwork_36_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_4_io_data_1_in_valid = PENetwork_16_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_4_io_data_1_in_bits = PENetwork_16_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_4_io_data_0_in_valid = PENetwork_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_4_io_data_0_in_bits = PENetwork_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_4_io_sig_stat2trans = _T_52_3; // @[pearray.scala 184:38]
  assign PE_5_clock = clock;
  assign PE_5_reset = reset;
  assign PE_5_io_data_2_in_valid = PENetwork_37_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_5_io_data_2_in_bits = PENetwork_37_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_5_io_data_1_in_valid = PENetwork_16_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_5_io_data_1_in_bits = PENetwork_16_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_5_io_data_0_in_valid = PENetwork_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_5_io_data_0_in_bits = PENetwork_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_5_io_sig_stat2trans = _T_62_3; // @[pearray.scala 184:38]
  assign PE_6_clock = clock;
  assign PE_6_reset = reset;
  assign PE_6_io_data_2_in_valid = PENetwork_38_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_6_io_data_2_in_bits = PENetwork_38_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_6_io_data_1_in_valid = PENetwork_16_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_6_io_data_1_in_bits = PENetwork_16_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_6_io_data_0_in_valid = PENetwork_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_6_io_data_0_in_bits = PENetwork_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_6_io_sig_stat2trans = _T_72_3; // @[pearray.scala 184:38]
  assign PE_7_clock = clock;
  assign PE_7_reset = reset;
  assign PE_7_io_data_2_in_valid = PENetwork_39_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_7_io_data_2_in_bits = PENetwork_39_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_7_io_data_1_in_valid = PENetwork_16_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_7_io_data_1_in_bits = PENetwork_16_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_7_io_data_0_in_valid = PENetwork_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_7_io_data_0_in_bits = PENetwork_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_7_io_sig_stat2trans = _T_82_3; // @[pearray.scala 184:38]
  assign PE_8_clock = clock;
  assign PE_8_reset = reset;
  assign PE_8_io_data_2_in_valid = PENetwork_40_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_8_io_data_2_in_bits = PENetwork_40_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_8_io_data_1_in_valid = PENetwork_16_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_8_io_data_1_in_bits = PENetwork_16_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_8_io_data_0_in_valid = PENetwork_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_8_io_data_0_in_bits = PENetwork_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_8_io_sig_stat2trans = _T_92_3; // @[pearray.scala 184:38]
  assign PE_9_clock = clock;
  assign PE_9_reset = reset;
  assign PE_9_io_data_2_in_valid = PENetwork_41_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_9_io_data_2_in_bits = PENetwork_41_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_9_io_data_1_in_valid = PENetwork_16_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_9_io_data_1_in_bits = PENetwork_16_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_9_io_data_0_in_valid = PENetwork_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_9_io_data_0_in_bits = PENetwork_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_9_io_sig_stat2trans = _T_102_3; // @[pearray.scala 184:38]
  assign PE_10_clock = clock;
  assign PE_10_reset = reset;
  assign PE_10_io_data_2_in_valid = PENetwork_42_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_10_io_data_2_in_bits = PENetwork_42_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_10_io_data_1_in_valid = PENetwork_16_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_10_io_data_1_in_bits = PENetwork_16_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_10_io_data_0_in_valid = PENetwork_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_10_io_data_0_in_bits = PENetwork_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_10_io_sig_stat2trans = _T_112_3; // @[pearray.scala 184:38]
  assign PE_11_clock = clock;
  assign PE_11_reset = reset;
  assign PE_11_io_data_2_in_valid = PENetwork_43_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_11_io_data_2_in_bits = PENetwork_43_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_11_io_data_1_in_valid = PENetwork_16_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_11_io_data_1_in_bits = PENetwork_16_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_11_io_data_0_in_valid = PENetwork_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_11_io_data_0_in_bits = PENetwork_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_11_io_sig_stat2trans = _T_122_3; // @[pearray.scala 184:38]
  assign PE_12_clock = clock;
  assign PE_12_reset = reset;
  assign PE_12_io_data_2_in_valid = PENetwork_44_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_12_io_data_2_in_bits = PENetwork_44_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_12_io_data_1_in_valid = PENetwork_16_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_12_io_data_1_in_bits = PENetwork_16_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_12_io_data_0_in_valid = PENetwork_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_12_io_data_0_in_bits = PENetwork_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_12_io_sig_stat2trans = _T_132_3; // @[pearray.scala 184:38]
  assign PE_13_clock = clock;
  assign PE_13_reset = reset;
  assign PE_13_io_data_2_in_valid = PENetwork_45_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_13_io_data_2_in_bits = PENetwork_45_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_13_io_data_1_in_valid = PENetwork_16_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_13_io_data_1_in_bits = PENetwork_16_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_13_io_data_0_in_valid = PENetwork_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_13_io_data_0_in_bits = PENetwork_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_13_io_sig_stat2trans = _T_142_3; // @[pearray.scala 184:38]
  assign PE_14_clock = clock;
  assign PE_14_reset = reset;
  assign PE_14_io_data_2_in_valid = PENetwork_46_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_14_io_data_2_in_bits = PENetwork_46_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_14_io_data_1_in_valid = PENetwork_16_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_14_io_data_1_in_bits = PENetwork_16_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_14_io_data_0_in_valid = PENetwork_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_14_io_data_0_in_bits = PENetwork_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_14_io_sig_stat2trans = _T_152_3; // @[pearray.scala 184:38]
  assign PE_15_clock = clock;
  assign PE_15_reset = reset;
  assign PE_15_io_data_2_in_valid = PENetwork_47_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_15_io_data_2_in_bits = PENetwork_47_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_15_io_data_1_in_valid = PENetwork_16_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_15_io_data_1_in_bits = PENetwork_16_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_15_io_data_0_in_valid = PENetwork_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_15_io_data_0_in_bits = PENetwork_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_15_io_sig_stat2trans = _T_162_3; // @[pearray.scala 184:38]
  assign PE_16_clock = clock;
  assign PE_16_reset = reset;
  assign PE_16_io_data_2_in_valid = PENetwork_32_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_16_io_data_2_in_bits = PENetwork_32_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_16_io_data_1_in_valid = PENetwork_17_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_16_io_data_1_in_bits = PENetwork_17_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_16_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_16_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_16_io_sig_stat2trans = _T_172_3; // @[pearray.scala 184:38]
  assign PE_17_clock = clock;
  assign PE_17_reset = reset;
  assign PE_17_io_data_2_in_valid = PENetwork_33_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_17_io_data_2_in_bits = PENetwork_33_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_17_io_data_1_in_valid = PENetwork_17_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_17_io_data_1_in_bits = PENetwork_17_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_17_io_data_0_in_valid = PENetwork_1_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_17_io_data_0_in_bits = PENetwork_1_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_17_io_sig_stat2trans = _T_182_3; // @[pearray.scala 184:38]
  assign PE_18_clock = clock;
  assign PE_18_reset = reset;
  assign PE_18_io_data_2_in_valid = PENetwork_34_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_18_io_data_2_in_bits = PENetwork_34_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_18_io_data_1_in_valid = PENetwork_17_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_18_io_data_1_in_bits = PENetwork_17_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_18_io_data_0_in_valid = PENetwork_1_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_18_io_data_0_in_bits = PENetwork_1_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_18_io_sig_stat2trans = _T_192_3; // @[pearray.scala 184:38]
  assign PE_19_clock = clock;
  assign PE_19_reset = reset;
  assign PE_19_io_data_2_in_valid = PENetwork_35_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_19_io_data_2_in_bits = PENetwork_35_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_19_io_data_1_in_valid = PENetwork_17_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_19_io_data_1_in_bits = PENetwork_17_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_19_io_data_0_in_valid = PENetwork_1_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_19_io_data_0_in_bits = PENetwork_1_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_19_io_sig_stat2trans = _T_202_3; // @[pearray.scala 184:38]
  assign PE_20_clock = clock;
  assign PE_20_reset = reset;
  assign PE_20_io_data_2_in_valid = PENetwork_36_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_20_io_data_2_in_bits = PENetwork_36_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_20_io_data_1_in_valid = PENetwork_17_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_20_io_data_1_in_bits = PENetwork_17_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_20_io_data_0_in_valid = PENetwork_1_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_20_io_data_0_in_bits = PENetwork_1_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_20_io_sig_stat2trans = _T_212_3; // @[pearray.scala 184:38]
  assign PE_21_clock = clock;
  assign PE_21_reset = reset;
  assign PE_21_io_data_2_in_valid = PENetwork_37_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_21_io_data_2_in_bits = PENetwork_37_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_21_io_data_1_in_valid = PENetwork_17_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_21_io_data_1_in_bits = PENetwork_17_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_21_io_data_0_in_valid = PENetwork_1_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_21_io_data_0_in_bits = PENetwork_1_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_21_io_sig_stat2trans = _T_222_3; // @[pearray.scala 184:38]
  assign PE_22_clock = clock;
  assign PE_22_reset = reset;
  assign PE_22_io_data_2_in_valid = PENetwork_38_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_22_io_data_2_in_bits = PENetwork_38_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_22_io_data_1_in_valid = PENetwork_17_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_22_io_data_1_in_bits = PENetwork_17_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_22_io_data_0_in_valid = PENetwork_1_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_22_io_data_0_in_bits = PENetwork_1_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_22_io_sig_stat2trans = _T_232_3; // @[pearray.scala 184:38]
  assign PE_23_clock = clock;
  assign PE_23_reset = reset;
  assign PE_23_io_data_2_in_valid = PENetwork_39_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_23_io_data_2_in_bits = PENetwork_39_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_23_io_data_1_in_valid = PENetwork_17_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_23_io_data_1_in_bits = PENetwork_17_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_23_io_data_0_in_valid = PENetwork_1_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_23_io_data_0_in_bits = PENetwork_1_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_23_io_sig_stat2trans = _T_242_3; // @[pearray.scala 184:38]
  assign PE_24_clock = clock;
  assign PE_24_reset = reset;
  assign PE_24_io_data_2_in_valid = PENetwork_40_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_24_io_data_2_in_bits = PENetwork_40_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_24_io_data_1_in_valid = PENetwork_17_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_24_io_data_1_in_bits = PENetwork_17_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_24_io_data_0_in_valid = PENetwork_1_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_24_io_data_0_in_bits = PENetwork_1_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_24_io_sig_stat2trans = _T_252_3; // @[pearray.scala 184:38]
  assign PE_25_clock = clock;
  assign PE_25_reset = reset;
  assign PE_25_io_data_2_in_valid = PENetwork_41_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_25_io_data_2_in_bits = PENetwork_41_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_25_io_data_1_in_valid = PENetwork_17_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_25_io_data_1_in_bits = PENetwork_17_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_25_io_data_0_in_valid = PENetwork_1_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_25_io_data_0_in_bits = PENetwork_1_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_25_io_sig_stat2trans = _T_262_3; // @[pearray.scala 184:38]
  assign PE_26_clock = clock;
  assign PE_26_reset = reset;
  assign PE_26_io_data_2_in_valid = PENetwork_42_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_26_io_data_2_in_bits = PENetwork_42_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_26_io_data_1_in_valid = PENetwork_17_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_26_io_data_1_in_bits = PENetwork_17_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_26_io_data_0_in_valid = PENetwork_1_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_26_io_data_0_in_bits = PENetwork_1_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_26_io_sig_stat2trans = _T_272_3; // @[pearray.scala 184:38]
  assign PE_27_clock = clock;
  assign PE_27_reset = reset;
  assign PE_27_io_data_2_in_valid = PENetwork_43_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_27_io_data_2_in_bits = PENetwork_43_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_27_io_data_1_in_valid = PENetwork_17_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_27_io_data_1_in_bits = PENetwork_17_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_27_io_data_0_in_valid = PENetwork_1_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_27_io_data_0_in_bits = PENetwork_1_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_27_io_sig_stat2trans = _T_282_3; // @[pearray.scala 184:38]
  assign PE_28_clock = clock;
  assign PE_28_reset = reset;
  assign PE_28_io_data_2_in_valid = PENetwork_44_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_28_io_data_2_in_bits = PENetwork_44_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_28_io_data_1_in_valid = PENetwork_17_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_28_io_data_1_in_bits = PENetwork_17_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_28_io_data_0_in_valid = PENetwork_1_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_28_io_data_0_in_bits = PENetwork_1_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_28_io_sig_stat2trans = _T_292_3; // @[pearray.scala 184:38]
  assign PE_29_clock = clock;
  assign PE_29_reset = reset;
  assign PE_29_io_data_2_in_valid = PENetwork_45_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_29_io_data_2_in_bits = PENetwork_45_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_29_io_data_1_in_valid = PENetwork_17_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_29_io_data_1_in_bits = PENetwork_17_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_29_io_data_0_in_valid = PENetwork_1_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_29_io_data_0_in_bits = PENetwork_1_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_29_io_sig_stat2trans = _T_302_3; // @[pearray.scala 184:38]
  assign PE_30_clock = clock;
  assign PE_30_reset = reset;
  assign PE_30_io_data_2_in_valid = PENetwork_46_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_30_io_data_2_in_bits = PENetwork_46_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_30_io_data_1_in_valid = PENetwork_17_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_30_io_data_1_in_bits = PENetwork_17_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_30_io_data_0_in_valid = PENetwork_1_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_30_io_data_0_in_bits = PENetwork_1_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_30_io_sig_stat2trans = _T_312_3; // @[pearray.scala 184:38]
  assign PE_31_clock = clock;
  assign PE_31_reset = reset;
  assign PE_31_io_data_2_in_valid = PENetwork_47_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_31_io_data_2_in_bits = PENetwork_47_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_31_io_data_1_in_valid = PENetwork_17_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_31_io_data_1_in_bits = PENetwork_17_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_31_io_data_0_in_valid = PENetwork_1_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_31_io_data_0_in_bits = PENetwork_1_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_31_io_sig_stat2trans = _T_322_3; // @[pearray.scala 184:38]
  assign PE_32_clock = clock;
  assign PE_32_reset = reset;
  assign PE_32_io_data_2_in_valid = PENetwork_32_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_32_io_data_2_in_bits = PENetwork_32_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_32_io_data_1_in_valid = PENetwork_18_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_32_io_data_1_in_bits = PENetwork_18_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_32_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_32_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_32_io_sig_stat2trans = _T_332_3; // @[pearray.scala 184:38]
  assign PE_33_clock = clock;
  assign PE_33_reset = reset;
  assign PE_33_io_data_2_in_valid = PENetwork_33_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_33_io_data_2_in_bits = PENetwork_33_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_33_io_data_1_in_valid = PENetwork_18_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_33_io_data_1_in_bits = PENetwork_18_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_33_io_data_0_in_valid = PENetwork_2_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_33_io_data_0_in_bits = PENetwork_2_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_33_io_sig_stat2trans = _T_342_3; // @[pearray.scala 184:38]
  assign PE_34_clock = clock;
  assign PE_34_reset = reset;
  assign PE_34_io_data_2_in_valid = PENetwork_34_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_34_io_data_2_in_bits = PENetwork_34_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_34_io_data_1_in_valid = PENetwork_18_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_34_io_data_1_in_bits = PENetwork_18_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_34_io_data_0_in_valid = PENetwork_2_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_34_io_data_0_in_bits = PENetwork_2_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_34_io_sig_stat2trans = _T_352_3; // @[pearray.scala 184:38]
  assign PE_35_clock = clock;
  assign PE_35_reset = reset;
  assign PE_35_io_data_2_in_valid = PENetwork_35_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_35_io_data_2_in_bits = PENetwork_35_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_35_io_data_1_in_valid = PENetwork_18_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_35_io_data_1_in_bits = PENetwork_18_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_35_io_data_0_in_valid = PENetwork_2_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_35_io_data_0_in_bits = PENetwork_2_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_35_io_sig_stat2trans = _T_362_3; // @[pearray.scala 184:38]
  assign PE_36_clock = clock;
  assign PE_36_reset = reset;
  assign PE_36_io_data_2_in_valid = PENetwork_36_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_36_io_data_2_in_bits = PENetwork_36_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_36_io_data_1_in_valid = PENetwork_18_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_36_io_data_1_in_bits = PENetwork_18_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_36_io_data_0_in_valid = PENetwork_2_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_36_io_data_0_in_bits = PENetwork_2_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_36_io_sig_stat2trans = _T_372_3; // @[pearray.scala 184:38]
  assign PE_37_clock = clock;
  assign PE_37_reset = reset;
  assign PE_37_io_data_2_in_valid = PENetwork_37_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_37_io_data_2_in_bits = PENetwork_37_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_37_io_data_1_in_valid = PENetwork_18_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_37_io_data_1_in_bits = PENetwork_18_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_37_io_data_0_in_valid = PENetwork_2_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_37_io_data_0_in_bits = PENetwork_2_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_37_io_sig_stat2trans = _T_382_3; // @[pearray.scala 184:38]
  assign PE_38_clock = clock;
  assign PE_38_reset = reset;
  assign PE_38_io_data_2_in_valid = PENetwork_38_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_38_io_data_2_in_bits = PENetwork_38_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_38_io_data_1_in_valid = PENetwork_18_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_38_io_data_1_in_bits = PENetwork_18_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_38_io_data_0_in_valid = PENetwork_2_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_38_io_data_0_in_bits = PENetwork_2_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_38_io_sig_stat2trans = _T_392_3; // @[pearray.scala 184:38]
  assign PE_39_clock = clock;
  assign PE_39_reset = reset;
  assign PE_39_io_data_2_in_valid = PENetwork_39_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_39_io_data_2_in_bits = PENetwork_39_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_39_io_data_1_in_valid = PENetwork_18_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_39_io_data_1_in_bits = PENetwork_18_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_39_io_data_0_in_valid = PENetwork_2_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_39_io_data_0_in_bits = PENetwork_2_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_39_io_sig_stat2trans = _T_402_3; // @[pearray.scala 184:38]
  assign PE_40_clock = clock;
  assign PE_40_reset = reset;
  assign PE_40_io_data_2_in_valid = PENetwork_40_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_40_io_data_2_in_bits = PENetwork_40_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_40_io_data_1_in_valid = PENetwork_18_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_40_io_data_1_in_bits = PENetwork_18_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_40_io_data_0_in_valid = PENetwork_2_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_40_io_data_0_in_bits = PENetwork_2_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_40_io_sig_stat2trans = _T_412_3; // @[pearray.scala 184:38]
  assign PE_41_clock = clock;
  assign PE_41_reset = reset;
  assign PE_41_io_data_2_in_valid = PENetwork_41_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_41_io_data_2_in_bits = PENetwork_41_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_41_io_data_1_in_valid = PENetwork_18_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_41_io_data_1_in_bits = PENetwork_18_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_41_io_data_0_in_valid = PENetwork_2_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_41_io_data_0_in_bits = PENetwork_2_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_41_io_sig_stat2trans = _T_422_3; // @[pearray.scala 184:38]
  assign PE_42_clock = clock;
  assign PE_42_reset = reset;
  assign PE_42_io_data_2_in_valid = PENetwork_42_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_42_io_data_2_in_bits = PENetwork_42_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_42_io_data_1_in_valid = PENetwork_18_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_42_io_data_1_in_bits = PENetwork_18_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_42_io_data_0_in_valid = PENetwork_2_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_42_io_data_0_in_bits = PENetwork_2_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_42_io_sig_stat2trans = _T_432_3; // @[pearray.scala 184:38]
  assign PE_43_clock = clock;
  assign PE_43_reset = reset;
  assign PE_43_io_data_2_in_valid = PENetwork_43_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_43_io_data_2_in_bits = PENetwork_43_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_43_io_data_1_in_valid = PENetwork_18_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_43_io_data_1_in_bits = PENetwork_18_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_43_io_data_0_in_valid = PENetwork_2_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_43_io_data_0_in_bits = PENetwork_2_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_43_io_sig_stat2trans = _T_442_3; // @[pearray.scala 184:38]
  assign PE_44_clock = clock;
  assign PE_44_reset = reset;
  assign PE_44_io_data_2_in_valid = PENetwork_44_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_44_io_data_2_in_bits = PENetwork_44_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_44_io_data_1_in_valid = PENetwork_18_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_44_io_data_1_in_bits = PENetwork_18_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_44_io_data_0_in_valid = PENetwork_2_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_44_io_data_0_in_bits = PENetwork_2_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_44_io_sig_stat2trans = _T_452_3; // @[pearray.scala 184:38]
  assign PE_45_clock = clock;
  assign PE_45_reset = reset;
  assign PE_45_io_data_2_in_valid = PENetwork_45_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_45_io_data_2_in_bits = PENetwork_45_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_45_io_data_1_in_valid = PENetwork_18_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_45_io_data_1_in_bits = PENetwork_18_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_45_io_data_0_in_valid = PENetwork_2_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_45_io_data_0_in_bits = PENetwork_2_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_45_io_sig_stat2trans = _T_462_3; // @[pearray.scala 184:38]
  assign PE_46_clock = clock;
  assign PE_46_reset = reset;
  assign PE_46_io_data_2_in_valid = PENetwork_46_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_46_io_data_2_in_bits = PENetwork_46_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_46_io_data_1_in_valid = PENetwork_18_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_46_io_data_1_in_bits = PENetwork_18_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_46_io_data_0_in_valid = PENetwork_2_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_46_io_data_0_in_bits = PENetwork_2_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_46_io_sig_stat2trans = _T_472_3; // @[pearray.scala 184:38]
  assign PE_47_clock = clock;
  assign PE_47_reset = reset;
  assign PE_47_io_data_2_in_valid = PENetwork_47_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_47_io_data_2_in_bits = PENetwork_47_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_47_io_data_1_in_valid = PENetwork_18_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_47_io_data_1_in_bits = PENetwork_18_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_47_io_data_0_in_valid = PENetwork_2_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_47_io_data_0_in_bits = PENetwork_2_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_47_io_sig_stat2trans = _T_482_3; // @[pearray.scala 184:38]
  assign PE_48_clock = clock;
  assign PE_48_reset = reset;
  assign PE_48_io_data_2_in_valid = PENetwork_32_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_48_io_data_2_in_bits = PENetwork_32_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_48_io_data_1_in_valid = PENetwork_19_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_48_io_data_1_in_bits = PENetwork_19_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_48_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_48_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_48_io_sig_stat2trans = _T_492_3; // @[pearray.scala 184:38]
  assign PE_49_clock = clock;
  assign PE_49_reset = reset;
  assign PE_49_io_data_2_in_valid = PENetwork_33_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_49_io_data_2_in_bits = PENetwork_33_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_49_io_data_1_in_valid = PENetwork_19_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_49_io_data_1_in_bits = PENetwork_19_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_49_io_data_0_in_valid = PENetwork_3_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_49_io_data_0_in_bits = PENetwork_3_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_49_io_sig_stat2trans = _T_502_3; // @[pearray.scala 184:38]
  assign PE_50_clock = clock;
  assign PE_50_reset = reset;
  assign PE_50_io_data_2_in_valid = PENetwork_34_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_50_io_data_2_in_bits = PENetwork_34_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_50_io_data_1_in_valid = PENetwork_19_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_50_io_data_1_in_bits = PENetwork_19_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_50_io_data_0_in_valid = PENetwork_3_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_50_io_data_0_in_bits = PENetwork_3_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_50_io_sig_stat2trans = _T_512_3; // @[pearray.scala 184:38]
  assign PE_51_clock = clock;
  assign PE_51_reset = reset;
  assign PE_51_io_data_2_in_valid = PENetwork_35_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_51_io_data_2_in_bits = PENetwork_35_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_51_io_data_1_in_valid = PENetwork_19_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_51_io_data_1_in_bits = PENetwork_19_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_51_io_data_0_in_valid = PENetwork_3_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_51_io_data_0_in_bits = PENetwork_3_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_51_io_sig_stat2trans = _T_522_3; // @[pearray.scala 184:38]
  assign PE_52_clock = clock;
  assign PE_52_reset = reset;
  assign PE_52_io_data_2_in_valid = PENetwork_36_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_52_io_data_2_in_bits = PENetwork_36_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_52_io_data_1_in_valid = PENetwork_19_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_52_io_data_1_in_bits = PENetwork_19_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_52_io_data_0_in_valid = PENetwork_3_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_52_io_data_0_in_bits = PENetwork_3_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_52_io_sig_stat2trans = _T_532_3; // @[pearray.scala 184:38]
  assign PE_53_clock = clock;
  assign PE_53_reset = reset;
  assign PE_53_io_data_2_in_valid = PENetwork_37_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_53_io_data_2_in_bits = PENetwork_37_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_53_io_data_1_in_valid = PENetwork_19_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_53_io_data_1_in_bits = PENetwork_19_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_53_io_data_0_in_valid = PENetwork_3_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_53_io_data_0_in_bits = PENetwork_3_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_53_io_sig_stat2trans = _T_542_3; // @[pearray.scala 184:38]
  assign PE_54_clock = clock;
  assign PE_54_reset = reset;
  assign PE_54_io_data_2_in_valid = PENetwork_38_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_54_io_data_2_in_bits = PENetwork_38_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_54_io_data_1_in_valid = PENetwork_19_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_54_io_data_1_in_bits = PENetwork_19_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_54_io_data_0_in_valid = PENetwork_3_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_54_io_data_0_in_bits = PENetwork_3_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_54_io_sig_stat2trans = _T_552_3; // @[pearray.scala 184:38]
  assign PE_55_clock = clock;
  assign PE_55_reset = reset;
  assign PE_55_io_data_2_in_valid = PENetwork_39_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_55_io_data_2_in_bits = PENetwork_39_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_55_io_data_1_in_valid = PENetwork_19_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_55_io_data_1_in_bits = PENetwork_19_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_55_io_data_0_in_valid = PENetwork_3_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_55_io_data_0_in_bits = PENetwork_3_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_55_io_sig_stat2trans = _T_562_3; // @[pearray.scala 184:38]
  assign PE_56_clock = clock;
  assign PE_56_reset = reset;
  assign PE_56_io_data_2_in_valid = PENetwork_40_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_56_io_data_2_in_bits = PENetwork_40_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_56_io_data_1_in_valid = PENetwork_19_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_56_io_data_1_in_bits = PENetwork_19_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_56_io_data_0_in_valid = PENetwork_3_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_56_io_data_0_in_bits = PENetwork_3_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_56_io_sig_stat2trans = _T_572_3; // @[pearray.scala 184:38]
  assign PE_57_clock = clock;
  assign PE_57_reset = reset;
  assign PE_57_io_data_2_in_valid = PENetwork_41_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_57_io_data_2_in_bits = PENetwork_41_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_57_io_data_1_in_valid = PENetwork_19_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_57_io_data_1_in_bits = PENetwork_19_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_57_io_data_0_in_valid = PENetwork_3_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_57_io_data_0_in_bits = PENetwork_3_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_57_io_sig_stat2trans = _T_582_3; // @[pearray.scala 184:38]
  assign PE_58_clock = clock;
  assign PE_58_reset = reset;
  assign PE_58_io_data_2_in_valid = PENetwork_42_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_58_io_data_2_in_bits = PENetwork_42_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_58_io_data_1_in_valid = PENetwork_19_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_58_io_data_1_in_bits = PENetwork_19_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_58_io_data_0_in_valid = PENetwork_3_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_58_io_data_0_in_bits = PENetwork_3_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_58_io_sig_stat2trans = _T_592_3; // @[pearray.scala 184:38]
  assign PE_59_clock = clock;
  assign PE_59_reset = reset;
  assign PE_59_io_data_2_in_valid = PENetwork_43_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_59_io_data_2_in_bits = PENetwork_43_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_59_io_data_1_in_valid = PENetwork_19_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_59_io_data_1_in_bits = PENetwork_19_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_59_io_data_0_in_valid = PENetwork_3_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_59_io_data_0_in_bits = PENetwork_3_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_59_io_sig_stat2trans = _T_602_3; // @[pearray.scala 184:38]
  assign PE_60_clock = clock;
  assign PE_60_reset = reset;
  assign PE_60_io_data_2_in_valid = PENetwork_44_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_60_io_data_2_in_bits = PENetwork_44_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_60_io_data_1_in_valid = PENetwork_19_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_60_io_data_1_in_bits = PENetwork_19_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_60_io_data_0_in_valid = PENetwork_3_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_60_io_data_0_in_bits = PENetwork_3_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_60_io_sig_stat2trans = _T_612_3; // @[pearray.scala 184:38]
  assign PE_61_clock = clock;
  assign PE_61_reset = reset;
  assign PE_61_io_data_2_in_valid = PENetwork_45_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_61_io_data_2_in_bits = PENetwork_45_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_61_io_data_1_in_valid = PENetwork_19_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_61_io_data_1_in_bits = PENetwork_19_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_61_io_data_0_in_valid = PENetwork_3_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_61_io_data_0_in_bits = PENetwork_3_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_61_io_sig_stat2trans = _T_622_3; // @[pearray.scala 184:38]
  assign PE_62_clock = clock;
  assign PE_62_reset = reset;
  assign PE_62_io_data_2_in_valid = PENetwork_46_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_62_io_data_2_in_bits = PENetwork_46_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_62_io_data_1_in_valid = PENetwork_19_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_62_io_data_1_in_bits = PENetwork_19_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_62_io_data_0_in_valid = PENetwork_3_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_62_io_data_0_in_bits = PENetwork_3_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_62_io_sig_stat2trans = _T_632_3; // @[pearray.scala 184:38]
  assign PE_63_clock = clock;
  assign PE_63_reset = reset;
  assign PE_63_io_data_2_in_valid = PENetwork_47_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_63_io_data_2_in_bits = PENetwork_47_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_63_io_data_1_in_valid = PENetwork_19_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_63_io_data_1_in_bits = PENetwork_19_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_63_io_data_0_in_valid = PENetwork_3_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_63_io_data_0_in_bits = PENetwork_3_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_63_io_sig_stat2trans = _T_642_3; // @[pearray.scala 184:38]
  assign PE_64_clock = clock;
  assign PE_64_reset = reset;
  assign PE_64_io_data_2_in_valid = PENetwork_32_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_64_io_data_2_in_bits = PENetwork_32_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_64_io_data_1_in_valid = PENetwork_20_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_64_io_data_1_in_bits = PENetwork_20_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_64_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_64_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_64_io_sig_stat2trans = _T_652_3; // @[pearray.scala 184:38]
  assign PE_65_clock = clock;
  assign PE_65_reset = reset;
  assign PE_65_io_data_2_in_valid = PENetwork_33_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_65_io_data_2_in_bits = PENetwork_33_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_65_io_data_1_in_valid = PENetwork_20_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_65_io_data_1_in_bits = PENetwork_20_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_65_io_data_0_in_valid = PENetwork_4_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_65_io_data_0_in_bits = PENetwork_4_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_65_io_sig_stat2trans = _T_662_3; // @[pearray.scala 184:38]
  assign PE_66_clock = clock;
  assign PE_66_reset = reset;
  assign PE_66_io_data_2_in_valid = PENetwork_34_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_66_io_data_2_in_bits = PENetwork_34_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_66_io_data_1_in_valid = PENetwork_20_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_66_io_data_1_in_bits = PENetwork_20_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_66_io_data_0_in_valid = PENetwork_4_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_66_io_data_0_in_bits = PENetwork_4_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_66_io_sig_stat2trans = _T_672_3; // @[pearray.scala 184:38]
  assign PE_67_clock = clock;
  assign PE_67_reset = reset;
  assign PE_67_io_data_2_in_valid = PENetwork_35_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_67_io_data_2_in_bits = PENetwork_35_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_67_io_data_1_in_valid = PENetwork_20_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_67_io_data_1_in_bits = PENetwork_20_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_67_io_data_0_in_valid = PENetwork_4_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_67_io_data_0_in_bits = PENetwork_4_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_67_io_sig_stat2trans = _T_682_3; // @[pearray.scala 184:38]
  assign PE_68_clock = clock;
  assign PE_68_reset = reset;
  assign PE_68_io_data_2_in_valid = PENetwork_36_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_68_io_data_2_in_bits = PENetwork_36_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_68_io_data_1_in_valid = PENetwork_20_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_68_io_data_1_in_bits = PENetwork_20_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_68_io_data_0_in_valid = PENetwork_4_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_68_io_data_0_in_bits = PENetwork_4_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_68_io_sig_stat2trans = _T_692_3; // @[pearray.scala 184:38]
  assign PE_69_clock = clock;
  assign PE_69_reset = reset;
  assign PE_69_io_data_2_in_valid = PENetwork_37_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_69_io_data_2_in_bits = PENetwork_37_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_69_io_data_1_in_valid = PENetwork_20_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_69_io_data_1_in_bits = PENetwork_20_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_69_io_data_0_in_valid = PENetwork_4_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_69_io_data_0_in_bits = PENetwork_4_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_69_io_sig_stat2trans = _T_702_3; // @[pearray.scala 184:38]
  assign PE_70_clock = clock;
  assign PE_70_reset = reset;
  assign PE_70_io_data_2_in_valid = PENetwork_38_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_70_io_data_2_in_bits = PENetwork_38_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_70_io_data_1_in_valid = PENetwork_20_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_70_io_data_1_in_bits = PENetwork_20_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_70_io_data_0_in_valid = PENetwork_4_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_70_io_data_0_in_bits = PENetwork_4_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_70_io_sig_stat2trans = _T_712_3; // @[pearray.scala 184:38]
  assign PE_71_clock = clock;
  assign PE_71_reset = reset;
  assign PE_71_io_data_2_in_valid = PENetwork_39_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_71_io_data_2_in_bits = PENetwork_39_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_71_io_data_1_in_valid = PENetwork_20_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_71_io_data_1_in_bits = PENetwork_20_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_71_io_data_0_in_valid = PENetwork_4_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_71_io_data_0_in_bits = PENetwork_4_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_71_io_sig_stat2trans = _T_722_3; // @[pearray.scala 184:38]
  assign PE_72_clock = clock;
  assign PE_72_reset = reset;
  assign PE_72_io_data_2_in_valid = PENetwork_40_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_72_io_data_2_in_bits = PENetwork_40_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_72_io_data_1_in_valid = PENetwork_20_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_72_io_data_1_in_bits = PENetwork_20_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_72_io_data_0_in_valid = PENetwork_4_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_72_io_data_0_in_bits = PENetwork_4_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_72_io_sig_stat2trans = _T_732_3; // @[pearray.scala 184:38]
  assign PE_73_clock = clock;
  assign PE_73_reset = reset;
  assign PE_73_io_data_2_in_valid = PENetwork_41_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_73_io_data_2_in_bits = PENetwork_41_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_73_io_data_1_in_valid = PENetwork_20_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_73_io_data_1_in_bits = PENetwork_20_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_73_io_data_0_in_valid = PENetwork_4_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_73_io_data_0_in_bits = PENetwork_4_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_73_io_sig_stat2trans = _T_742_3; // @[pearray.scala 184:38]
  assign PE_74_clock = clock;
  assign PE_74_reset = reset;
  assign PE_74_io_data_2_in_valid = PENetwork_42_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_74_io_data_2_in_bits = PENetwork_42_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_74_io_data_1_in_valid = PENetwork_20_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_74_io_data_1_in_bits = PENetwork_20_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_74_io_data_0_in_valid = PENetwork_4_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_74_io_data_0_in_bits = PENetwork_4_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_74_io_sig_stat2trans = _T_752_3; // @[pearray.scala 184:38]
  assign PE_75_clock = clock;
  assign PE_75_reset = reset;
  assign PE_75_io_data_2_in_valid = PENetwork_43_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_75_io_data_2_in_bits = PENetwork_43_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_75_io_data_1_in_valid = PENetwork_20_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_75_io_data_1_in_bits = PENetwork_20_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_75_io_data_0_in_valid = PENetwork_4_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_75_io_data_0_in_bits = PENetwork_4_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_75_io_sig_stat2trans = _T_762_3; // @[pearray.scala 184:38]
  assign PE_76_clock = clock;
  assign PE_76_reset = reset;
  assign PE_76_io_data_2_in_valid = PENetwork_44_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_76_io_data_2_in_bits = PENetwork_44_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_76_io_data_1_in_valid = PENetwork_20_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_76_io_data_1_in_bits = PENetwork_20_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_76_io_data_0_in_valid = PENetwork_4_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_76_io_data_0_in_bits = PENetwork_4_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_76_io_sig_stat2trans = _T_772_3; // @[pearray.scala 184:38]
  assign PE_77_clock = clock;
  assign PE_77_reset = reset;
  assign PE_77_io_data_2_in_valid = PENetwork_45_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_77_io_data_2_in_bits = PENetwork_45_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_77_io_data_1_in_valid = PENetwork_20_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_77_io_data_1_in_bits = PENetwork_20_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_77_io_data_0_in_valid = PENetwork_4_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_77_io_data_0_in_bits = PENetwork_4_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_77_io_sig_stat2trans = _T_782_3; // @[pearray.scala 184:38]
  assign PE_78_clock = clock;
  assign PE_78_reset = reset;
  assign PE_78_io_data_2_in_valid = PENetwork_46_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_78_io_data_2_in_bits = PENetwork_46_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_78_io_data_1_in_valid = PENetwork_20_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_78_io_data_1_in_bits = PENetwork_20_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_78_io_data_0_in_valid = PENetwork_4_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_78_io_data_0_in_bits = PENetwork_4_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_78_io_sig_stat2trans = _T_792_3; // @[pearray.scala 184:38]
  assign PE_79_clock = clock;
  assign PE_79_reset = reset;
  assign PE_79_io_data_2_in_valid = PENetwork_47_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_79_io_data_2_in_bits = PENetwork_47_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_79_io_data_1_in_valid = PENetwork_20_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_79_io_data_1_in_bits = PENetwork_20_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_79_io_data_0_in_valid = PENetwork_4_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_79_io_data_0_in_bits = PENetwork_4_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_79_io_sig_stat2trans = _T_802_3; // @[pearray.scala 184:38]
  assign PE_80_clock = clock;
  assign PE_80_reset = reset;
  assign PE_80_io_data_2_in_valid = PENetwork_32_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_80_io_data_2_in_bits = PENetwork_32_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_80_io_data_1_in_valid = PENetwork_21_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_80_io_data_1_in_bits = PENetwork_21_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_80_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_80_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_80_io_sig_stat2trans = _T_812_3; // @[pearray.scala 184:38]
  assign PE_81_clock = clock;
  assign PE_81_reset = reset;
  assign PE_81_io_data_2_in_valid = PENetwork_33_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_81_io_data_2_in_bits = PENetwork_33_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_81_io_data_1_in_valid = PENetwork_21_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_81_io_data_1_in_bits = PENetwork_21_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_81_io_data_0_in_valid = PENetwork_5_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_81_io_data_0_in_bits = PENetwork_5_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_81_io_sig_stat2trans = _T_822_3; // @[pearray.scala 184:38]
  assign PE_82_clock = clock;
  assign PE_82_reset = reset;
  assign PE_82_io_data_2_in_valid = PENetwork_34_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_82_io_data_2_in_bits = PENetwork_34_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_82_io_data_1_in_valid = PENetwork_21_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_82_io_data_1_in_bits = PENetwork_21_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_82_io_data_0_in_valid = PENetwork_5_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_82_io_data_0_in_bits = PENetwork_5_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_82_io_sig_stat2trans = _T_832_3; // @[pearray.scala 184:38]
  assign PE_83_clock = clock;
  assign PE_83_reset = reset;
  assign PE_83_io_data_2_in_valid = PENetwork_35_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_83_io_data_2_in_bits = PENetwork_35_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_83_io_data_1_in_valid = PENetwork_21_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_83_io_data_1_in_bits = PENetwork_21_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_83_io_data_0_in_valid = PENetwork_5_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_83_io_data_0_in_bits = PENetwork_5_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_83_io_sig_stat2trans = _T_842_3; // @[pearray.scala 184:38]
  assign PE_84_clock = clock;
  assign PE_84_reset = reset;
  assign PE_84_io_data_2_in_valid = PENetwork_36_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_84_io_data_2_in_bits = PENetwork_36_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_84_io_data_1_in_valid = PENetwork_21_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_84_io_data_1_in_bits = PENetwork_21_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_84_io_data_0_in_valid = PENetwork_5_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_84_io_data_0_in_bits = PENetwork_5_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_84_io_sig_stat2trans = _T_852_3; // @[pearray.scala 184:38]
  assign PE_85_clock = clock;
  assign PE_85_reset = reset;
  assign PE_85_io_data_2_in_valid = PENetwork_37_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_85_io_data_2_in_bits = PENetwork_37_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_85_io_data_1_in_valid = PENetwork_21_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_85_io_data_1_in_bits = PENetwork_21_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_85_io_data_0_in_valid = PENetwork_5_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_85_io_data_0_in_bits = PENetwork_5_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_85_io_sig_stat2trans = _T_862_3; // @[pearray.scala 184:38]
  assign PE_86_clock = clock;
  assign PE_86_reset = reset;
  assign PE_86_io_data_2_in_valid = PENetwork_38_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_86_io_data_2_in_bits = PENetwork_38_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_86_io_data_1_in_valid = PENetwork_21_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_86_io_data_1_in_bits = PENetwork_21_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_86_io_data_0_in_valid = PENetwork_5_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_86_io_data_0_in_bits = PENetwork_5_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_86_io_sig_stat2trans = _T_872_3; // @[pearray.scala 184:38]
  assign PE_87_clock = clock;
  assign PE_87_reset = reset;
  assign PE_87_io_data_2_in_valid = PENetwork_39_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_87_io_data_2_in_bits = PENetwork_39_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_87_io_data_1_in_valid = PENetwork_21_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_87_io_data_1_in_bits = PENetwork_21_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_87_io_data_0_in_valid = PENetwork_5_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_87_io_data_0_in_bits = PENetwork_5_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_87_io_sig_stat2trans = _T_882_3; // @[pearray.scala 184:38]
  assign PE_88_clock = clock;
  assign PE_88_reset = reset;
  assign PE_88_io_data_2_in_valid = PENetwork_40_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_88_io_data_2_in_bits = PENetwork_40_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_88_io_data_1_in_valid = PENetwork_21_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_88_io_data_1_in_bits = PENetwork_21_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_88_io_data_0_in_valid = PENetwork_5_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_88_io_data_0_in_bits = PENetwork_5_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_88_io_sig_stat2trans = _T_892_3; // @[pearray.scala 184:38]
  assign PE_89_clock = clock;
  assign PE_89_reset = reset;
  assign PE_89_io_data_2_in_valid = PENetwork_41_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_89_io_data_2_in_bits = PENetwork_41_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_89_io_data_1_in_valid = PENetwork_21_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_89_io_data_1_in_bits = PENetwork_21_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_89_io_data_0_in_valid = PENetwork_5_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_89_io_data_0_in_bits = PENetwork_5_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_89_io_sig_stat2trans = _T_902_3; // @[pearray.scala 184:38]
  assign PE_90_clock = clock;
  assign PE_90_reset = reset;
  assign PE_90_io_data_2_in_valid = PENetwork_42_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_90_io_data_2_in_bits = PENetwork_42_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_90_io_data_1_in_valid = PENetwork_21_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_90_io_data_1_in_bits = PENetwork_21_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_90_io_data_0_in_valid = PENetwork_5_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_90_io_data_0_in_bits = PENetwork_5_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_90_io_sig_stat2trans = _T_912_3; // @[pearray.scala 184:38]
  assign PE_91_clock = clock;
  assign PE_91_reset = reset;
  assign PE_91_io_data_2_in_valid = PENetwork_43_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_91_io_data_2_in_bits = PENetwork_43_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_91_io_data_1_in_valid = PENetwork_21_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_91_io_data_1_in_bits = PENetwork_21_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_91_io_data_0_in_valid = PENetwork_5_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_91_io_data_0_in_bits = PENetwork_5_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_91_io_sig_stat2trans = _T_922_3; // @[pearray.scala 184:38]
  assign PE_92_clock = clock;
  assign PE_92_reset = reset;
  assign PE_92_io_data_2_in_valid = PENetwork_44_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_92_io_data_2_in_bits = PENetwork_44_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_92_io_data_1_in_valid = PENetwork_21_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_92_io_data_1_in_bits = PENetwork_21_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_92_io_data_0_in_valid = PENetwork_5_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_92_io_data_0_in_bits = PENetwork_5_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_92_io_sig_stat2trans = _T_932_3; // @[pearray.scala 184:38]
  assign PE_93_clock = clock;
  assign PE_93_reset = reset;
  assign PE_93_io_data_2_in_valid = PENetwork_45_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_93_io_data_2_in_bits = PENetwork_45_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_93_io_data_1_in_valid = PENetwork_21_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_93_io_data_1_in_bits = PENetwork_21_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_93_io_data_0_in_valid = PENetwork_5_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_93_io_data_0_in_bits = PENetwork_5_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_93_io_sig_stat2trans = _T_942_3; // @[pearray.scala 184:38]
  assign PE_94_clock = clock;
  assign PE_94_reset = reset;
  assign PE_94_io_data_2_in_valid = PENetwork_46_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_94_io_data_2_in_bits = PENetwork_46_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_94_io_data_1_in_valid = PENetwork_21_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_94_io_data_1_in_bits = PENetwork_21_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_94_io_data_0_in_valid = PENetwork_5_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_94_io_data_0_in_bits = PENetwork_5_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_94_io_sig_stat2trans = _T_952_3; // @[pearray.scala 184:38]
  assign PE_95_clock = clock;
  assign PE_95_reset = reset;
  assign PE_95_io_data_2_in_valid = PENetwork_47_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_95_io_data_2_in_bits = PENetwork_47_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_95_io_data_1_in_valid = PENetwork_21_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_95_io_data_1_in_bits = PENetwork_21_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_95_io_data_0_in_valid = PENetwork_5_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_95_io_data_0_in_bits = PENetwork_5_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_95_io_sig_stat2trans = _T_962_3; // @[pearray.scala 184:38]
  assign PE_96_clock = clock;
  assign PE_96_reset = reset;
  assign PE_96_io_data_2_in_valid = PENetwork_32_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_96_io_data_2_in_bits = PENetwork_32_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_96_io_data_1_in_valid = PENetwork_22_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_96_io_data_1_in_bits = PENetwork_22_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_96_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_96_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_96_io_sig_stat2trans = _T_972_3; // @[pearray.scala 184:38]
  assign PE_97_clock = clock;
  assign PE_97_reset = reset;
  assign PE_97_io_data_2_in_valid = PENetwork_33_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_97_io_data_2_in_bits = PENetwork_33_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_97_io_data_1_in_valid = PENetwork_22_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_97_io_data_1_in_bits = PENetwork_22_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_97_io_data_0_in_valid = PENetwork_6_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_97_io_data_0_in_bits = PENetwork_6_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_97_io_sig_stat2trans = _T_982_3; // @[pearray.scala 184:38]
  assign PE_98_clock = clock;
  assign PE_98_reset = reset;
  assign PE_98_io_data_2_in_valid = PENetwork_34_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_98_io_data_2_in_bits = PENetwork_34_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_98_io_data_1_in_valid = PENetwork_22_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_98_io_data_1_in_bits = PENetwork_22_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_98_io_data_0_in_valid = PENetwork_6_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_98_io_data_0_in_bits = PENetwork_6_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_98_io_sig_stat2trans = _T_992_3; // @[pearray.scala 184:38]
  assign PE_99_clock = clock;
  assign PE_99_reset = reset;
  assign PE_99_io_data_2_in_valid = PENetwork_35_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_99_io_data_2_in_bits = PENetwork_35_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_99_io_data_1_in_valid = PENetwork_22_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_99_io_data_1_in_bits = PENetwork_22_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_99_io_data_0_in_valid = PENetwork_6_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_99_io_data_0_in_bits = PENetwork_6_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_99_io_sig_stat2trans = _T_1002_3; // @[pearray.scala 184:38]
  assign PE_100_clock = clock;
  assign PE_100_reset = reset;
  assign PE_100_io_data_2_in_valid = PENetwork_36_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_100_io_data_2_in_bits = PENetwork_36_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_100_io_data_1_in_valid = PENetwork_22_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_100_io_data_1_in_bits = PENetwork_22_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_100_io_data_0_in_valid = PENetwork_6_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_100_io_data_0_in_bits = PENetwork_6_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_100_io_sig_stat2trans = _T_1012_3; // @[pearray.scala 184:38]
  assign PE_101_clock = clock;
  assign PE_101_reset = reset;
  assign PE_101_io_data_2_in_valid = PENetwork_37_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_101_io_data_2_in_bits = PENetwork_37_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_101_io_data_1_in_valid = PENetwork_22_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_101_io_data_1_in_bits = PENetwork_22_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_101_io_data_0_in_valid = PENetwork_6_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_101_io_data_0_in_bits = PENetwork_6_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_101_io_sig_stat2trans = _T_1022_3; // @[pearray.scala 184:38]
  assign PE_102_clock = clock;
  assign PE_102_reset = reset;
  assign PE_102_io_data_2_in_valid = PENetwork_38_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_102_io_data_2_in_bits = PENetwork_38_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_102_io_data_1_in_valid = PENetwork_22_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_102_io_data_1_in_bits = PENetwork_22_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_102_io_data_0_in_valid = PENetwork_6_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_102_io_data_0_in_bits = PENetwork_6_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_102_io_sig_stat2trans = _T_1032_3; // @[pearray.scala 184:38]
  assign PE_103_clock = clock;
  assign PE_103_reset = reset;
  assign PE_103_io_data_2_in_valid = PENetwork_39_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_103_io_data_2_in_bits = PENetwork_39_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_103_io_data_1_in_valid = PENetwork_22_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_103_io_data_1_in_bits = PENetwork_22_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_103_io_data_0_in_valid = PENetwork_6_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_103_io_data_0_in_bits = PENetwork_6_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_103_io_sig_stat2trans = _T_1042_3; // @[pearray.scala 184:38]
  assign PE_104_clock = clock;
  assign PE_104_reset = reset;
  assign PE_104_io_data_2_in_valid = PENetwork_40_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_104_io_data_2_in_bits = PENetwork_40_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_104_io_data_1_in_valid = PENetwork_22_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_104_io_data_1_in_bits = PENetwork_22_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_104_io_data_0_in_valid = PENetwork_6_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_104_io_data_0_in_bits = PENetwork_6_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_104_io_sig_stat2trans = _T_1052_3; // @[pearray.scala 184:38]
  assign PE_105_clock = clock;
  assign PE_105_reset = reset;
  assign PE_105_io_data_2_in_valid = PENetwork_41_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_105_io_data_2_in_bits = PENetwork_41_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_105_io_data_1_in_valid = PENetwork_22_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_105_io_data_1_in_bits = PENetwork_22_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_105_io_data_0_in_valid = PENetwork_6_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_105_io_data_0_in_bits = PENetwork_6_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_105_io_sig_stat2trans = _T_1062_3; // @[pearray.scala 184:38]
  assign PE_106_clock = clock;
  assign PE_106_reset = reset;
  assign PE_106_io_data_2_in_valid = PENetwork_42_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_106_io_data_2_in_bits = PENetwork_42_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_106_io_data_1_in_valid = PENetwork_22_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_106_io_data_1_in_bits = PENetwork_22_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_106_io_data_0_in_valid = PENetwork_6_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_106_io_data_0_in_bits = PENetwork_6_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_106_io_sig_stat2trans = _T_1072_3; // @[pearray.scala 184:38]
  assign PE_107_clock = clock;
  assign PE_107_reset = reset;
  assign PE_107_io_data_2_in_valid = PENetwork_43_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_107_io_data_2_in_bits = PENetwork_43_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_107_io_data_1_in_valid = PENetwork_22_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_107_io_data_1_in_bits = PENetwork_22_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_107_io_data_0_in_valid = PENetwork_6_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_107_io_data_0_in_bits = PENetwork_6_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_107_io_sig_stat2trans = _T_1082_3; // @[pearray.scala 184:38]
  assign PE_108_clock = clock;
  assign PE_108_reset = reset;
  assign PE_108_io_data_2_in_valid = PENetwork_44_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_108_io_data_2_in_bits = PENetwork_44_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_108_io_data_1_in_valid = PENetwork_22_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_108_io_data_1_in_bits = PENetwork_22_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_108_io_data_0_in_valid = PENetwork_6_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_108_io_data_0_in_bits = PENetwork_6_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_108_io_sig_stat2trans = _T_1092_3; // @[pearray.scala 184:38]
  assign PE_109_clock = clock;
  assign PE_109_reset = reset;
  assign PE_109_io_data_2_in_valid = PENetwork_45_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_109_io_data_2_in_bits = PENetwork_45_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_109_io_data_1_in_valid = PENetwork_22_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_109_io_data_1_in_bits = PENetwork_22_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_109_io_data_0_in_valid = PENetwork_6_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_109_io_data_0_in_bits = PENetwork_6_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_109_io_sig_stat2trans = _T_1102_3; // @[pearray.scala 184:38]
  assign PE_110_clock = clock;
  assign PE_110_reset = reset;
  assign PE_110_io_data_2_in_valid = PENetwork_46_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_110_io_data_2_in_bits = PENetwork_46_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_110_io_data_1_in_valid = PENetwork_22_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_110_io_data_1_in_bits = PENetwork_22_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_110_io_data_0_in_valid = PENetwork_6_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_110_io_data_0_in_bits = PENetwork_6_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_110_io_sig_stat2trans = _T_1112_3; // @[pearray.scala 184:38]
  assign PE_111_clock = clock;
  assign PE_111_reset = reset;
  assign PE_111_io_data_2_in_valid = PENetwork_47_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_111_io_data_2_in_bits = PENetwork_47_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_111_io_data_1_in_valid = PENetwork_22_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_111_io_data_1_in_bits = PENetwork_22_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_111_io_data_0_in_valid = PENetwork_6_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_111_io_data_0_in_bits = PENetwork_6_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_111_io_sig_stat2trans = _T_1122_3; // @[pearray.scala 184:38]
  assign PE_112_clock = clock;
  assign PE_112_reset = reset;
  assign PE_112_io_data_2_in_valid = PENetwork_32_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_112_io_data_2_in_bits = PENetwork_32_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_112_io_data_1_in_valid = PENetwork_23_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_112_io_data_1_in_bits = PENetwork_23_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_112_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_112_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_112_io_sig_stat2trans = _T_1132_3; // @[pearray.scala 184:38]
  assign PE_113_clock = clock;
  assign PE_113_reset = reset;
  assign PE_113_io_data_2_in_valid = PENetwork_33_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_113_io_data_2_in_bits = PENetwork_33_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_113_io_data_1_in_valid = PENetwork_23_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_113_io_data_1_in_bits = PENetwork_23_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_113_io_data_0_in_valid = PENetwork_7_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_113_io_data_0_in_bits = PENetwork_7_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_113_io_sig_stat2trans = _T_1142_3; // @[pearray.scala 184:38]
  assign PE_114_clock = clock;
  assign PE_114_reset = reset;
  assign PE_114_io_data_2_in_valid = PENetwork_34_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_114_io_data_2_in_bits = PENetwork_34_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_114_io_data_1_in_valid = PENetwork_23_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_114_io_data_1_in_bits = PENetwork_23_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_114_io_data_0_in_valid = PENetwork_7_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_114_io_data_0_in_bits = PENetwork_7_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_114_io_sig_stat2trans = _T_1152_3; // @[pearray.scala 184:38]
  assign PE_115_clock = clock;
  assign PE_115_reset = reset;
  assign PE_115_io_data_2_in_valid = PENetwork_35_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_115_io_data_2_in_bits = PENetwork_35_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_115_io_data_1_in_valid = PENetwork_23_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_115_io_data_1_in_bits = PENetwork_23_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_115_io_data_0_in_valid = PENetwork_7_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_115_io_data_0_in_bits = PENetwork_7_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_115_io_sig_stat2trans = _T_1162_3; // @[pearray.scala 184:38]
  assign PE_116_clock = clock;
  assign PE_116_reset = reset;
  assign PE_116_io_data_2_in_valid = PENetwork_36_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_116_io_data_2_in_bits = PENetwork_36_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_116_io_data_1_in_valid = PENetwork_23_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_116_io_data_1_in_bits = PENetwork_23_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_116_io_data_0_in_valid = PENetwork_7_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_116_io_data_0_in_bits = PENetwork_7_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_116_io_sig_stat2trans = _T_1172_3; // @[pearray.scala 184:38]
  assign PE_117_clock = clock;
  assign PE_117_reset = reset;
  assign PE_117_io_data_2_in_valid = PENetwork_37_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_117_io_data_2_in_bits = PENetwork_37_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_117_io_data_1_in_valid = PENetwork_23_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_117_io_data_1_in_bits = PENetwork_23_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_117_io_data_0_in_valid = PENetwork_7_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_117_io_data_0_in_bits = PENetwork_7_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_117_io_sig_stat2trans = _T_1182_3; // @[pearray.scala 184:38]
  assign PE_118_clock = clock;
  assign PE_118_reset = reset;
  assign PE_118_io_data_2_in_valid = PENetwork_38_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_118_io_data_2_in_bits = PENetwork_38_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_118_io_data_1_in_valid = PENetwork_23_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_118_io_data_1_in_bits = PENetwork_23_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_118_io_data_0_in_valid = PENetwork_7_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_118_io_data_0_in_bits = PENetwork_7_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_118_io_sig_stat2trans = _T_1192_3; // @[pearray.scala 184:38]
  assign PE_119_clock = clock;
  assign PE_119_reset = reset;
  assign PE_119_io_data_2_in_valid = PENetwork_39_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_119_io_data_2_in_bits = PENetwork_39_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_119_io_data_1_in_valid = PENetwork_23_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_119_io_data_1_in_bits = PENetwork_23_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_119_io_data_0_in_valid = PENetwork_7_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_119_io_data_0_in_bits = PENetwork_7_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_119_io_sig_stat2trans = _T_1202_3; // @[pearray.scala 184:38]
  assign PE_120_clock = clock;
  assign PE_120_reset = reset;
  assign PE_120_io_data_2_in_valid = PENetwork_40_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_120_io_data_2_in_bits = PENetwork_40_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_120_io_data_1_in_valid = PENetwork_23_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_120_io_data_1_in_bits = PENetwork_23_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_120_io_data_0_in_valid = PENetwork_7_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_120_io_data_0_in_bits = PENetwork_7_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_120_io_sig_stat2trans = _T_1212_3; // @[pearray.scala 184:38]
  assign PE_121_clock = clock;
  assign PE_121_reset = reset;
  assign PE_121_io_data_2_in_valid = PENetwork_41_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_121_io_data_2_in_bits = PENetwork_41_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_121_io_data_1_in_valid = PENetwork_23_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_121_io_data_1_in_bits = PENetwork_23_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_121_io_data_0_in_valid = PENetwork_7_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_121_io_data_0_in_bits = PENetwork_7_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_121_io_sig_stat2trans = _T_1222_3; // @[pearray.scala 184:38]
  assign PE_122_clock = clock;
  assign PE_122_reset = reset;
  assign PE_122_io_data_2_in_valid = PENetwork_42_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_122_io_data_2_in_bits = PENetwork_42_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_122_io_data_1_in_valid = PENetwork_23_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_122_io_data_1_in_bits = PENetwork_23_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_122_io_data_0_in_valid = PENetwork_7_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_122_io_data_0_in_bits = PENetwork_7_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_122_io_sig_stat2trans = _T_1232_3; // @[pearray.scala 184:38]
  assign PE_123_clock = clock;
  assign PE_123_reset = reset;
  assign PE_123_io_data_2_in_valid = PENetwork_43_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_123_io_data_2_in_bits = PENetwork_43_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_123_io_data_1_in_valid = PENetwork_23_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_123_io_data_1_in_bits = PENetwork_23_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_123_io_data_0_in_valid = PENetwork_7_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_123_io_data_0_in_bits = PENetwork_7_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_123_io_sig_stat2trans = _T_1242_3; // @[pearray.scala 184:38]
  assign PE_124_clock = clock;
  assign PE_124_reset = reset;
  assign PE_124_io_data_2_in_valid = PENetwork_44_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_124_io_data_2_in_bits = PENetwork_44_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_124_io_data_1_in_valid = PENetwork_23_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_124_io_data_1_in_bits = PENetwork_23_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_124_io_data_0_in_valid = PENetwork_7_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_124_io_data_0_in_bits = PENetwork_7_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_124_io_sig_stat2trans = _T_1252_3; // @[pearray.scala 184:38]
  assign PE_125_clock = clock;
  assign PE_125_reset = reset;
  assign PE_125_io_data_2_in_valid = PENetwork_45_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_125_io_data_2_in_bits = PENetwork_45_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_125_io_data_1_in_valid = PENetwork_23_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_125_io_data_1_in_bits = PENetwork_23_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_125_io_data_0_in_valid = PENetwork_7_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_125_io_data_0_in_bits = PENetwork_7_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_125_io_sig_stat2trans = _T_1262_3; // @[pearray.scala 184:38]
  assign PE_126_clock = clock;
  assign PE_126_reset = reset;
  assign PE_126_io_data_2_in_valid = PENetwork_46_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_126_io_data_2_in_bits = PENetwork_46_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_126_io_data_1_in_valid = PENetwork_23_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_126_io_data_1_in_bits = PENetwork_23_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_126_io_data_0_in_valid = PENetwork_7_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_126_io_data_0_in_bits = PENetwork_7_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_126_io_sig_stat2trans = _T_1272_3; // @[pearray.scala 184:38]
  assign PE_127_clock = clock;
  assign PE_127_reset = reset;
  assign PE_127_io_data_2_in_valid = PENetwork_47_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_127_io_data_2_in_bits = PENetwork_47_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_127_io_data_1_in_valid = PENetwork_23_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_127_io_data_1_in_bits = PENetwork_23_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_127_io_data_0_in_valid = PENetwork_7_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_127_io_data_0_in_bits = PENetwork_7_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_127_io_sig_stat2trans = _T_1282_3; // @[pearray.scala 184:38]
  assign PE_128_clock = clock;
  assign PE_128_reset = reset;
  assign PE_128_io_data_2_in_valid = PENetwork_32_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_128_io_data_2_in_bits = PENetwork_32_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_128_io_data_1_in_valid = PENetwork_24_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_128_io_data_1_in_bits = PENetwork_24_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_128_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_128_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_128_io_sig_stat2trans = _T_1292_3; // @[pearray.scala 184:38]
  assign PE_129_clock = clock;
  assign PE_129_reset = reset;
  assign PE_129_io_data_2_in_valid = PENetwork_33_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_129_io_data_2_in_bits = PENetwork_33_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_129_io_data_1_in_valid = PENetwork_24_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_129_io_data_1_in_bits = PENetwork_24_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_129_io_data_0_in_valid = PENetwork_8_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_129_io_data_0_in_bits = PENetwork_8_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_129_io_sig_stat2trans = _T_1302_3; // @[pearray.scala 184:38]
  assign PE_130_clock = clock;
  assign PE_130_reset = reset;
  assign PE_130_io_data_2_in_valid = PENetwork_34_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_130_io_data_2_in_bits = PENetwork_34_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_130_io_data_1_in_valid = PENetwork_24_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_130_io_data_1_in_bits = PENetwork_24_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_130_io_data_0_in_valid = PENetwork_8_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_130_io_data_0_in_bits = PENetwork_8_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_130_io_sig_stat2trans = _T_1312_3; // @[pearray.scala 184:38]
  assign PE_131_clock = clock;
  assign PE_131_reset = reset;
  assign PE_131_io_data_2_in_valid = PENetwork_35_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_131_io_data_2_in_bits = PENetwork_35_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_131_io_data_1_in_valid = PENetwork_24_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_131_io_data_1_in_bits = PENetwork_24_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_131_io_data_0_in_valid = PENetwork_8_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_131_io_data_0_in_bits = PENetwork_8_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_131_io_sig_stat2trans = _T_1322_3; // @[pearray.scala 184:38]
  assign PE_132_clock = clock;
  assign PE_132_reset = reset;
  assign PE_132_io_data_2_in_valid = PENetwork_36_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_132_io_data_2_in_bits = PENetwork_36_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_132_io_data_1_in_valid = PENetwork_24_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_132_io_data_1_in_bits = PENetwork_24_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_132_io_data_0_in_valid = PENetwork_8_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_132_io_data_0_in_bits = PENetwork_8_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_132_io_sig_stat2trans = _T_1332_3; // @[pearray.scala 184:38]
  assign PE_133_clock = clock;
  assign PE_133_reset = reset;
  assign PE_133_io_data_2_in_valid = PENetwork_37_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_133_io_data_2_in_bits = PENetwork_37_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_133_io_data_1_in_valid = PENetwork_24_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_133_io_data_1_in_bits = PENetwork_24_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_133_io_data_0_in_valid = PENetwork_8_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_133_io_data_0_in_bits = PENetwork_8_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_133_io_sig_stat2trans = _T_1342_3; // @[pearray.scala 184:38]
  assign PE_134_clock = clock;
  assign PE_134_reset = reset;
  assign PE_134_io_data_2_in_valid = PENetwork_38_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_134_io_data_2_in_bits = PENetwork_38_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_134_io_data_1_in_valid = PENetwork_24_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_134_io_data_1_in_bits = PENetwork_24_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_134_io_data_0_in_valid = PENetwork_8_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_134_io_data_0_in_bits = PENetwork_8_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_134_io_sig_stat2trans = _T_1352_3; // @[pearray.scala 184:38]
  assign PE_135_clock = clock;
  assign PE_135_reset = reset;
  assign PE_135_io_data_2_in_valid = PENetwork_39_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_135_io_data_2_in_bits = PENetwork_39_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_135_io_data_1_in_valid = PENetwork_24_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_135_io_data_1_in_bits = PENetwork_24_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_135_io_data_0_in_valid = PENetwork_8_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_135_io_data_0_in_bits = PENetwork_8_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_135_io_sig_stat2trans = _T_1362_3; // @[pearray.scala 184:38]
  assign PE_136_clock = clock;
  assign PE_136_reset = reset;
  assign PE_136_io_data_2_in_valid = PENetwork_40_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_136_io_data_2_in_bits = PENetwork_40_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_136_io_data_1_in_valid = PENetwork_24_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_136_io_data_1_in_bits = PENetwork_24_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_136_io_data_0_in_valid = PENetwork_8_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_136_io_data_0_in_bits = PENetwork_8_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_136_io_sig_stat2trans = _T_1372_3; // @[pearray.scala 184:38]
  assign PE_137_clock = clock;
  assign PE_137_reset = reset;
  assign PE_137_io_data_2_in_valid = PENetwork_41_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_137_io_data_2_in_bits = PENetwork_41_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_137_io_data_1_in_valid = PENetwork_24_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_137_io_data_1_in_bits = PENetwork_24_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_137_io_data_0_in_valid = PENetwork_8_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_137_io_data_0_in_bits = PENetwork_8_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_137_io_sig_stat2trans = _T_1382_3; // @[pearray.scala 184:38]
  assign PE_138_clock = clock;
  assign PE_138_reset = reset;
  assign PE_138_io_data_2_in_valid = PENetwork_42_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_138_io_data_2_in_bits = PENetwork_42_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_138_io_data_1_in_valid = PENetwork_24_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_138_io_data_1_in_bits = PENetwork_24_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_138_io_data_0_in_valid = PENetwork_8_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_138_io_data_0_in_bits = PENetwork_8_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_138_io_sig_stat2trans = _T_1392_3; // @[pearray.scala 184:38]
  assign PE_139_clock = clock;
  assign PE_139_reset = reset;
  assign PE_139_io_data_2_in_valid = PENetwork_43_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_139_io_data_2_in_bits = PENetwork_43_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_139_io_data_1_in_valid = PENetwork_24_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_139_io_data_1_in_bits = PENetwork_24_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_139_io_data_0_in_valid = PENetwork_8_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_139_io_data_0_in_bits = PENetwork_8_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_139_io_sig_stat2trans = _T_1402_3; // @[pearray.scala 184:38]
  assign PE_140_clock = clock;
  assign PE_140_reset = reset;
  assign PE_140_io_data_2_in_valid = PENetwork_44_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_140_io_data_2_in_bits = PENetwork_44_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_140_io_data_1_in_valid = PENetwork_24_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_140_io_data_1_in_bits = PENetwork_24_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_140_io_data_0_in_valid = PENetwork_8_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_140_io_data_0_in_bits = PENetwork_8_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_140_io_sig_stat2trans = _T_1412_3; // @[pearray.scala 184:38]
  assign PE_141_clock = clock;
  assign PE_141_reset = reset;
  assign PE_141_io_data_2_in_valid = PENetwork_45_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_141_io_data_2_in_bits = PENetwork_45_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_141_io_data_1_in_valid = PENetwork_24_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_141_io_data_1_in_bits = PENetwork_24_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_141_io_data_0_in_valid = PENetwork_8_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_141_io_data_0_in_bits = PENetwork_8_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_141_io_sig_stat2trans = _T_1422_3; // @[pearray.scala 184:38]
  assign PE_142_clock = clock;
  assign PE_142_reset = reset;
  assign PE_142_io_data_2_in_valid = PENetwork_46_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_142_io_data_2_in_bits = PENetwork_46_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_142_io_data_1_in_valid = PENetwork_24_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_142_io_data_1_in_bits = PENetwork_24_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_142_io_data_0_in_valid = PENetwork_8_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_142_io_data_0_in_bits = PENetwork_8_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_142_io_sig_stat2trans = _T_1432_3; // @[pearray.scala 184:38]
  assign PE_143_clock = clock;
  assign PE_143_reset = reset;
  assign PE_143_io_data_2_in_valid = PENetwork_47_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_143_io_data_2_in_bits = PENetwork_47_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_143_io_data_1_in_valid = PENetwork_24_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_143_io_data_1_in_bits = PENetwork_24_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_143_io_data_0_in_valid = PENetwork_8_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_143_io_data_0_in_bits = PENetwork_8_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_143_io_sig_stat2trans = _T_1442_3; // @[pearray.scala 184:38]
  assign PE_144_clock = clock;
  assign PE_144_reset = reset;
  assign PE_144_io_data_2_in_valid = PENetwork_32_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_144_io_data_2_in_bits = PENetwork_32_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_144_io_data_1_in_valid = PENetwork_25_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_144_io_data_1_in_bits = PENetwork_25_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_144_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_144_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_144_io_sig_stat2trans = _T_1452_3; // @[pearray.scala 184:38]
  assign PE_145_clock = clock;
  assign PE_145_reset = reset;
  assign PE_145_io_data_2_in_valid = PENetwork_33_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_145_io_data_2_in_bits = PENetwork_33_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_145_io_data_1_in_valid = PENetwork_25_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_145_io_data_1_in_bits = PENetwork_25_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_145_io_data_0_in_valid = PENetwork_9_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_145_io_data_0_in_bits = PENetwork_9_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_145_io_sig_stat2trans = _T_1462_3; // @[pearray.scala 184:38]
  assign PE_146_clock = clock;
  assign PE_146_reset = reset;
  assign PE_146_io_data_2_in_valid = PENetwork_34_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_146_io_data_2_in_bits = PENetwork_34_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_146_io_data_1_in_valid = PENetwork_25_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_146_io_data_1_in_bits = PENetwork_25_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_146_io_data_0_in_valid = PENetwork_9_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_146_io_data_0_in_bits = PENetwork_9_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_146_io_sig_stat2trans = _T_1472_3; // @[pearray.scala 184:38]
  assign PE_147_clock = clock;
  assign PE_147_reset = reset;
  assign PE_147_io_data_2_in_valid = PENetwork_35_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_147_io_data_2_in_bits = PENetwork_35_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_147_io_data_1_in_valid = PENetwork_25_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_147_io_data_1_in_bits = PENetwork_25_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_147_io_data_0_in_valid = PENetwork_9_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_147_io_data_0_in_bits = PENetwork_9_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_147_io_sig_stat2trans = _T_1482_3; // @[pearray.scala 184:38]
  assign PE_148_clock = clock;
  assign PE_148_reset = reset;
  assign PE_148_io_data_2_in_valid = PENetwork_36_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_148_io_data_2_in_bits = PENetwork_36_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_148_io_data_1_in_valid = PENetwork_25_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_148_io_data_1_in_bits = PENetwork_25_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_148_io_data_0_in_valid = PENetwork_9_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_148_io_data_0_in_bits = PENetwork_9_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_148_io_sig_stat2trans = _T_1492_3; // @[pearray.scala 184:38]
  assign PE_149_clock = clock;
  assign PE_149_reset = reset;
  assign PE_149_io_data_2_in_valid = PENetwork_37_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_149_io_data_2_in_bits = PENetwork_37_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_149_io_data_1_in_valid = PENetwork_25_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_149_io_data_1_in_bits = PENetwork_25_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_149_io_data_0_in_valid = PENetwork_9_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_149_io_data_0_in_bits = PENetwork_9_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_149_io_sig_stat2trans = _T_1502_3; // @[pearray.scala 184:38]
  assign PE_150_clock = clock;
  assign PE_150_reset = reset;
  assign PE_150_io_data_2_in_valid = PENetwork_38_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_150_io_data_2_in_bits = PENetwork_38_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_150_io_data_1_in_valid = PENetwork_25_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_150_io_data_1_in_bits = PENetwork_25_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_150_io_data_0_in_valid = PENetwork_9_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_150_io_data_0_in_bits = PENetwork_9_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_150_io_sig_stat2trans = _T_1512_3; // @[pearray.scala 184:38]
  assign PE_151_clock = clock;
  assign PE_151_reset = reset;
  assign PE_151_io_data_2_in_valid = PENetwork_39_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_151_io_data_2_in_bits = PENetwork_39_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_151_io_data_1_in_valid = PENetwork_25_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_151_io_data_1_in_bits = PENetwork_25_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_151_io_data_0_in_valid = PENetwork_9_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_151_io_data_0_in_bits = PENetwork_9_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_151_io_sig_stat2trans = _T_1522_3; // @[pearray.scala 184:38]
  assign PE_152_clock = clock;
  assign PE_152_reset = reset;
  assign PE_152_io_data_2_in_valid = PENetwork_40_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_152_io_data_2_in_bits = PENetwork_40_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_152_io_data_1_in_valid = PENetwork_25_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_152_io_data_1_in_bits = PENetwork_25_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_152_io_data_0_in_valid = PENetwork_9_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_152_io_data_0_in_bits = PENetwork_9_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_152_io_sig_stat2trans = _T_1532_3; // @[pearray.scala 184:38]
  assign PE_153_clock = clock;
  assign PE_153_reset = reset;
  assign PE_153_io_data_2_in_valid = PENetwork_41_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_153_io_data_2_in_bits = PENetwork_41_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_153_io_data_1_in_valid = PENetwork_25_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_153_io_data_1_in_bits = PENetwork_25_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_153_io_data_0_in_valid = PENetwork_9_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_153_io_data_0_in_bits = PENetwork_9_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_153_io_sig_stat2trans = _T_1542_3; // @[pearray.scala 184:38]
  assign PE_154_clock = clock;
  assign PE_154_reset = reset;
  assign PE_154_io_data_2_in_valid = PENetwork_42_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_154_io_data_2_in_bits = PENetwork_42_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_154_io_data_1_in_valid = PENetwork_25_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_154_io_data_1_in_bits = PENetwork_25_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_154_io_data_0_in_valid = PENetwork_9_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_154_io_data_0_in_bits = PENetwork_9_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_154_io_sig_stat2trans = _T_1552_3; // @[pearray.scala 184:38]
  assign PE_155_clock = clock;
  assign PE_155_reset = reset;
  assign PE_155_io_data_2_in_valid = PENetwork_43_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_155_io_data_2_in_bits = PENetwork_43_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_155_io_data_1_in_valid = PENetwork_25_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_155_io_data_1_in_bits = PENetwork_25_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_155_io_data_0_in_valid = PENetwork_9_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_155_io_data_0_in_bits = PENetwork_9_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_155_io_sig_stat2trans = _T_1562_3; // @[pearray.scala 184:38]
  assign PE_156_clock = clock;
  assign PE_156_reset = reset;
  assign PE_156_io_data_2_in_valid = PENetwork_44_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_156_io_data_2_in_bits = PENetwork_44_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_156_io_data_1_in_valid = PENetwork_25_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_156_io_data_1_in_bits = PENetwork_25_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_156_io_data_0_in_valid = PENetwork_9_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_156_io_data_0_in_bits = PENetwork_9_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_156_io_sig_stat2trans = _T_1572_3; // @[pearray.scala 184:38]
  assign PE_157_clock = clock;
  assign PE_157_reset = reset;
  assign PE_157_io_data_2_in_valid = PENetwork_45_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_157_io_data_2_in_bits = PENetwork_45_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_157_io_data_1_in_valid = PENetwork_25_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_157_io_data_1_in_bits = PENetwork_25_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_157_io_data_0_in_valid = PENetwork_9_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_157_io_data_0_in_bits = PENetwork_9_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_157_io_sig_stat2trans = _T_1582_3; // @[pearray.scala 184:38]
  assign PE_158_clock = clock;
  assign PE_158_reset = reset;
  assign PE_158_io_data_2_in_valid = PENetwork_46_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_158_io_data_2_in_bits = PENetwork_46_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_158_io_data_1_in_valid = PENetwork_25_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_158_io_data_1_in_bits = PENetwork_25_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_158_io_data_0_in_valid = PENetwork_9_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_158_io_data_0_in_bits = PENetwork_9_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_158_io_sig_stat2trans = _T_1592_3; // @[pearray.scala 184:38]
  assign PE_159_clock = clock;
  assign PE_159_reset = reset;
  assign PE_159_io_data_2_in_valid = PENetwork_47_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_159_io_data_2_in_bits = PENetwork_47_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_159_io_data_1_in_valid = PENetwork_25_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_159_io_data_1_in_bits = PENetwork_25_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_159_io_data_0_in_valid = PENetwork_9_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_159_io_data_0_in_bits = PENetwork_9_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_159_io_sig_stat2trans = _T_1602_3; // @[pearray.scala 184:38]
  assign PE_160_clock = clock;
  assign PE_160_reset = reset;
  assign PE_160_io_data_2_in_valid = PENetwork_32_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_160_io_data_2_in_bits = PENetwork_32_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_160_io_data_1_in_valid = PENetwork_26_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_160_io_data_1_in_bits = PENetwork_26_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_160_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_160_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_160_io_sig_stat2trans = _T_1612_3; // @[pearray.scala 184:38]
  assign PE_161_clock = clock;
  assign PE_161_reset = reset;
  assign PE_161_io_data_2_in_valid = PENetwork_33_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_161_io_data_2_in_bits = PENetwork_33_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_161_io_data_1_in_valid = PENetwork_26_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_161_io_data_1_in_bits = PENetwork_26_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_161_io_data_0_in_valid = PENetwork_10_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_161_io_data_0_in_bits = PENetwork_10_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_161_io_sig_stat2trans = _T_1622_3; // @[pearray.scala 184:38]
  assign PE_162_clock = clock;
  assign PE_162_reset = reset;
  assign PE_162_io_data_2_in_valid = PENetwork_34_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_162_io_data_2_in_bits = PENetwork_34_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_162_io_data_1_in_valid = PENetwork_26_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_162_io_data_1_in_bits = PENetwork_26_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_162_io_data_0_in_valid = PENetwork_10_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_162_io_data_0_in_bits = PENetwork_10_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_162_io_sig_stat2trans = _T_1632_3; // @[pearray.scala 184:38]
  assign PE_163_clock = clock;
  assign PE_163_reset = reset;
  assign PE_163_io_data_2_in_valid = PENetwork_35_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_163_io_data_2_in_bits = PENetwork_35_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_163_io_data_1_in_valid = PENetwork_26_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_163_io_data_1_in_bits = PENetwork_26_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_163_io_data_0_in_valid = PENetwork_10_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_163_io_data_0_in_bits = PENetwork_10_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_163_io_sig_stat2trans = _T_1642_3; // @[pearray.scala 184:38]
  assign PE_164_clock = clock;
  assign PE_164_reset = reset;
  assign PE_164_io_data_2_in_valid = PENetwork_36_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_164_io_data_2_in_bits = PENetwork_36_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_164_io_data_1_in_valid = PENetwork_26_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_164_io_data_1_in_bits = PENetwork_26_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_164_io_data_0_in_valid = PENetwork_10_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_164_io_data_0_in_bits = PENetwork_10_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_164_io_sig_stat2trans = _T_1652_3; // @[pearray.scala 184:38]
  assign PE_165_clock = clock;
  assign PE_165_reset = reset;
  assign PE_165_io_data_2_in_valid = PENetwork_37_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_165_io_data_2_in_bits = PENetwork_37_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_165_io_data_1_in_valid = PENetwork_26_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_165_io_data_1_in_bits = PENetwork_26_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_165_io_data_0_in_valid = PENetwork_10_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_165_io_data_0_in_bits = PENetwork_10_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_165_io_sig_stat2trans = _T_1662_3; // @[pearray.scala 184:38]
  assign PE_166_clock = clock;
  assign PE_166_reset = reset;
  assign PE_166_io_data_2_in_valid = PENetwork_38_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_166_io_data_2_in_bits = PENetwork_38_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_166_io_data_1_in_valid = PENetwork_26_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_166_io_data_1_in_bits = PENetwork_26_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_166_io_data_0_in_valid = PENetwork_10_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_166_io_data_0_in_bits = PENetwork_10_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_166_io_sig_stat2trans = _T_1672_3; // @[pearray.scala 184:38]
  assign PE_167_clock = clock;
  assign PE_167_reset = reset;
  assign PE_167_io_data_2_in_valid = PENetwork_39_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_167_io_data_2_in_bits = PENetwork_39_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_167_io_data_1_in_valid = PENetwork_26_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_167_io_data_1_in_bits = PENetwork_26_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_167_io_data_0_in_valid = PENetwork_10_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_167_io_data_0_in_bits = PENetwork_10_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_167_io_sig_stat2trans = _T_1682_3; // @[pearray.scala 184:38]
  assign PE_168_clock = clock;
  assign PE_168_reset = reset;
  assign PE_168_io_data_2_in_valid = PENetwork_40_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_168_io_data_2_in_bits = PENetwork_40_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_168_io_data_1_in_valid = PENetwork_26_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_168_io_data_1_in_bits = PENetwork_26_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_168_io_data_0_in_valid = PENetwork_10_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_168_io_data_0_in_bits = PENetwork_10_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_168_io_sig_stat2trans = _T_1692_3; // @[pearray.scala 184:38]
  assign PE_169_clock = clock;
  assign PE_169_reset = reset;
  assign PE_169_io_data_2_in_valid = PENetwork_41_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_169_io_data_2_in_bits = PENetwork_41_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_169_io_data_1_in_valid = PENetwork_26_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_169_io_data_1_in_bits = PENetwork_26_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_169_io_data_0_in_valid = PENetwork_10_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_169_io_data_0_in_bits = PENetwork_10_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_169_io_sig_stat2trans = _T_1702_3; // @[pearray.scala 184:38]
  assign PE_170_clock = clock;
  assign PE_170_reset = reset;
  assign PE_170_io_data_2_in_valid = PENetwork_42_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_170_io_data_2_in_bits = PENetwork_42_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_170_io_data_1_in_valid = PENetwork_26_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_170_io_data_1_in_bits = PENetwork_26_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_170_io_data_0_in_valid = PENetwork_10_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_170_io_data_0_in_bits = PENetwork_10_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_170_io_sig_stat2trans = _T_1712_3; // @[pearray.scala 184:38]
  assign PE_171_clock = clock;
  assign PE_171_reset = reset;
  assign PE_171_io_data_2_in_valid = PENetwork_43_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_171_io_data_2_in_bits = PENetwork_43_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_171_io_data_1_in_valid = PENetwork_26_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_171_io_data_1_in_bits = PENetwork_26_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_171_io_data_0_in_valid = PENetwork_10_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_171_io_data_0_in_bits = PENetwork_10_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_171_io_sig_stat2trans = _T_1722_3; // @[pearray.scala 184:38]
  assign PE_172_clock = clock;
  assign PE_172_reset = reset;
  assign PE_172_io_data_2_in_valid = PENetwork_44_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_172_io_data_2_in_bits = PENetwork_44_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_172_io_data_1_in_valid = PENetwork_26_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_172_io_data_1_in_bits = PENetwork_26_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_172_io_data_0_in_valid = PENetwork_10_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_172_io_data_0_in_bits = PENetwork_10_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_172_io_sig_stat2trans = _T_1732_3; // @[pearray.scala 184:38]
  assign PE_173_clock = clock;
  assign PE_173_reset = reset;
  assign PE_173_io_data_2_in_valid = PENetwork_45_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_173_io_data_2_in_bits = PENetwork_45_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_173_io_data_1_in_valid = PENetwork_26_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_173_io_data_1_in_bits = PENetwork_26_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_173_io_data_0_in_valid = PENetwork_10_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_173_io_data_0_in_bits = PENetwork_10_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_173_io_sig_stat2trans = _T_1742_3; // @[pearray.scala 184:38]
  assign PE_174_clock = clock;
  assign PE_174_reset = reset;
  assign PE_174_io_data_2_in_valid = PENetwork_46_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_174_io_data_2_in_bits = PENetwork_46_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_174_io_data_1_in_valid = PENetwork_26_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_174_io_data_1_in_bits = PENetwork_26_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_174_io_data_0_in_valid = PENetwork_10_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_174_io_data_0_in_bits = PENetwork_10_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_174_io_sig_stat2trans = _T_1752_3; // @[pearray.scala 184:38]
  assign PE_175_clock = clock;
  assign PE_175_reset = reset;
  assign PE_175_io_data_2_in_valid = PENetwork_47_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_175_io_data_2_in_bits = PENetwork_47_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_175_io_data_1_in_valid = PENetwork_26_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_175_io_data_1_in_bits = PENetwork_26_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_175_io_data_0_in_valid = PENetwork_10_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_175_io_data_0_in_bits = PENetwork_10_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_175_io_sig_stat2trans = _T_1762_3; // @[pearray.scala 184:38]
  assign PE_176_clock = clock;
  assign PE_176_reset = reset;
  assign PE_176_io_data_2_in_valid = PENetwork_32_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_176_io_data_2_in_bits = PENetwork_32_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_176_io_data_1_in_valid = PENetwork_27_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_176_io_data_1_in_bits = PENetwork_27_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_176_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_176_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_176_io_sig_stat2trans = _T_1772_3; // @[pearray.scala 184:38]
  assign PE_177_clock = clock;
  assign PE_177_reset = reset;
  assign PE_177_io_data_2_in_valid = PENetwork_33_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_177_io_data_2_in_bits = PENetwork_33_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_177_io_data_1_in_valid = PENetwork_27_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_177_io_data_1_in_bits = PENetwork_27_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_177_io_data_0_in_valid = PENetwork_11_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_177_io_data_0_in_bits = PENetwork_11_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_177_io_sig_stat2trans = _T_1782_3; // @[pearray.scala 184:38]
  assign PE_178_clock = clock;
  assign PE_178_reset = reset;
  assign PE_178_io_data_2_in_valid = PENetwork_34_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_178_io_data_2_in_bits = PENetwork_34_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_178_io_data_1_in_valid = PENetwork_27_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_178_io_data_1_in_bits = PENetwork_27_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_178_io_data_0_in_valid = PENetwork_11_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_178_io_data_0_in_bits = PENetwork_11_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_178_io_sig_stat2trans = _T_1792_3; // @[pearray.scala 184:38]
  assign PE_179_clock = clock;
  assign PE_179_reset = reset;
  assign PE_179_io_data_2_in_valid = PENetwork_35_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_179_io_data_2_in_bits = PENetwork_35_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_179_io_data_1_in_valid = PENetwork_27_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_179_io_data_1_in_bits = PENetwork_27_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_179_io_data_0_in_valid = PENetwork_11_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_179_io_data_0_in_bits = PENetwork_11_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_179_io_sig_stat2trans = _T_1802_3; // @[pearray.scala 184:38]
  assign PE_180_clock = clock;
  assign PE_180_reset = reset;
  assign PE_180_io_data_2_in_valid = PENetwork_36_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_180_io_data_2_in_bits = PENetwork_36_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_180_io_data_1_in_valid = PENetwork_27_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_180_io_data_1_in_bits = PENetwork_27_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_180_io_data_0_in_valid = PENetwork_11_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_180_io_data_0_in_bits = PENetwork_11_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_180_io_sig_stat2trans = _T_1812_3; // @[pearray.scala 184:38]
  assign PE_181_clock = clock;
  assign PE_181_reset = reset;
  assign PE_181_io_data_2_in_valid = PENetwork_37_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_181_io_data_2_in_bits = PENetwork_37_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_181_io_data_1_in_valid = PENetwork_27_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_181_io_data_1_in_bits = PENetwork_27_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_181_io_data_0_in_valid = PENetwork_11_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_181_io_data_0_in_bits = PENetwork_11_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_181_io_sig_stat2trans = _T_1822_3; // @[pearray.scala 184:38]
  assign PE_182_clock = clock;
  assign PE_182_reset = reset;
  assign PE_182_io_data_2_in_valid = PENetwork_38_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_182_io_data_2_in_bits = PENetwork_38_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_182_io_data_1_in_valid = PENetwork_27_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_182_io_data_1_in_bits = PENetwork_27_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_182_io_data_0_in_valid = PENetwork_11_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_182_io_data_0_in_bits = PENetwork_11_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_182_io_sig_stat2trans = _T_1832_3; // @[pearray.scala 184:38]
  assign PE_183_clock = clock;
  assign PE_183_reset = reset;
  assign PE_183_io_data_2_in_valid = PENetwork_39_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_183_io_data_2_in_bits = PENetwork_39_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_183_io_data_1_in_valid = PENetwork_27_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_183_io_data_1_in_bits = PENetwork_27_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_183_io_data_0_in_valid = PENetwork_11_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_183_io_data_0_in_bits = PENetwork_11_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_183_io_sig_stat2trans = _T_1842_3; // @[pearray.scala 184:38]
  assign PE_184_clock = clock;
  assign PE_184_reset = reset;
  assign PE_184_io_data_2_in_valid = PENetwork_40_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_184_io_data_2_in_bits = PENetwork_40_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_184_io_data_1_in_valid = PENetwork_27_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_184_io_data_1_in_bits = PENetwork_27_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_184_io_data_0_in_valid = PENetwork_11_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_184_io_data_0_in_bits = PENetwork_11_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_184_io_sig_stat2trans = _T_1852_3; // @[pearray.scala 184:38]
  assign PE_185_clock = clock;
  assign PE_185_reset = reset;
  assign PE_185_io_data_2_in_valid = PENetwork_41_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_185_io_data_2_in_bits = PENetwork_41_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_185_io_data_1_in_valid = PENetwork_27_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_185_io_data_1_in_bits = PENetwork_27_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_185_io_data_0_in_valid = PENetwork_11_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_185_io_data_0_in_bits = PENetwork_11_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_185_io_sig_stat2trans = _T_1862_3; // @[pearray.scala 184:38]
  assign PE_186_clock = clock;
  assign PE_186_reset = reset;
  assign PE_186_io_data_2_in_valid = PENetwork_42_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_186_io_data_2_in_bits = PENetwork_42_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_186_io_data_1_in_valid = PENetwork_27_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_186_io_data_1_in_bits = PENetwork_27_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_186_io_data_0_in_valid = PENetwork_11_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_186_io_data_0_in_bits = PENetwork_11_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_186_io_sig_stat2trans = _T_1872_3; // @[pearray.scala 184:38]
  assign PE_187_clock = clock;
  assign PE_187_reset = reset;
  assign PE_187_io_data_2_in_valid = PENetwork_43_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_187_io_data_2_in_bits = PENetwork_43_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_187_io_data_1_in_valid = PENetwork_27_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_187_io_data_1_in_bits = PENetwork_27_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_187_io_data_0_in_valid = PENetwork_11_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_187_io_data_0_in_bits = PENetwork_11_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_187_io_sig_stat2trans = _T_1882_3; // @[pearray.scala 184:38]
  assign PE_188_clock = clock;
  assign PE_188_reset = reset;
  assign PE_188_io_data_2_in_valid = PENetwork_44_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_188_io_data_2_in_bits = PENetwork_44_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_188_io_data_1_in_valid = PENetwork_27_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_188_io_data_1_in_bits = PENetwork_27_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_188_io_data_0_in_valid = PENetwork_11_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_188_io_data_0_in_bits = PENetwork_11_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_188_io_sig_stat2trans = _T_1892_3; // @[pearray.scala 184:38]
  assign PE_189_clock = clock;
  assign PE_189_reset = reset;
  assign PE_189_io_data_2_in_valid = PENetwork_45_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_189_io_data_2_in_bits = PENetwork_45_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_189_io_data_1_in_valid = PENetwork_27_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_189_io_data_1_in_bits = PENetwork_27_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_189_io_data_0_in_valid = PENetwork_11_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_189_io_data_0_in_bits = PENetwork_11_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_189_io_sig_stat2trans = _T_1902_3; // @[pearray.scala 184:38]
  assign PE_190_clock = clock;
  assign PE_190_reset = reset;
  assign PE_190_io_data_2_in_valid = PENetwork_46_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_190_io_data_2_in_bits = PENetwork_46_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_190_io_data_1_in_valid = PENetwork_27_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_190_io_data_1_in_bits = PENetwork_27_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_190_io_data_0_in_valid = PENetwork_11_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_190_io_data_0_in_bits = PENetwork_11_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_190_io_sig_stat2trans = _T_1912_3; // @[pearray.scala 184:38]
  assign PE_191_clock = clock;
  assign PE_191_reset = reset;
  assign PE_191_io_data_2_in_valid = PENetwork_47_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_191_io_data_2_in_bits = PENetwork_47_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_191_io_data_1_in_valid = PENetwork_27_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_191_io_data_1_in_bits = PENetwork_27_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_191_io_data_0_in_valid = PENetwork_11_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_191_io_data_0_in_bits = PENetwork_11_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_191_io_sig_stat2trans = _T_1922_3; // @[pearray.scala 184:38]
  assign PE_192_clock = clock;
  assign PE_192_reset = reset;
  assign PE_192_io_data_2_in_valid = PENetwork_32_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_192_io_data_2_in_bits = PENetwork_32_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_192_io_data_1_in_valid = PENetwork_28_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_192_io_data_1_in_bits = PENetwork_28_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_192_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_192_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_192_io_sig_stat2trans = _T_1932_3; // @[pearray.scala 184:38]
  assign PE_193_clock = clock;
  assign PE_193_reset = reset;
  assign PE_193_io_data_2_in_valid = PENetwork_33_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_193_io_data_2_in_bits = PENetwork_33_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_193_io_data_1_in_valid = PENetwork_28_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_193_io_data_1_in_bits = PENetwork_28_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_193_io_data_0_in_valid = PENetwork_12_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_193_io_data_0_in_bits = PENetwork_12_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_193_io_sig_stat2trans = _T_1942_3; // @[pearray.scala 184:38]
  assign PE_194_clock = clock;
  assign PE_194_reset = reset;
  assign PE_194_io_data_2_in_valid = PENetwork_34_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_194_io_data_2_in_bits = PENetwork_34_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_194_io_data_1_in_valid = PENetwork_28_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_194_io_data_1_in_bits = PENetwork_28_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_194_io_data_0_in_valid = PENetwork_12_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_194_io_data_0_in_bits = PENetwork_12_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_194_io_sig_stat2trans = _T_1952_3; // @[pearray.scala 184:38]
  assign PE_195_clock = clock;
  assign PE_195_reset = reset;
  assign PE_195_io_data_2_in_valid = PENetwork_35_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_195_io_data_2_in_bits = PENetwork_35_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_195_io_data_1_in_valid = PENetwork_28_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_195_io_data_1_in_bits = PENetwork_28_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_195_io_data_0_in_valid = PENetwork_12_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_195_io_data_0_in_bits = PENetwork_12_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_195_io_sig_stat2trans = _T_1962_3; // @[pearray.scala 184:38]
  assign PE_196_clock = clock;
  assign PE_196_reset = reset;
  assign PE_196_io_data_2_in_valid = PENetwork_36_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_196_io_data_2_in_bits = PENetwork_36_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_196_io_data_1_in_valid = PENetwork_28_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_196_io_data_1_in_bits = PENetwork_28_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_196_io_data_0_in_valid = PENetwork_12_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_196_io_data_0_in_bits = PENetwork_12_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_196_io_sig_stat2trans = _T_1972_3; // @[pearray.scala 184:38]
  assign PE_197_clock = clock;
  assign PE_197_reset = reset;
  assign PE_197_io_data_2_in_valid = PENetwork_37_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_197_io_data_2_in_bits = PENetwork_37_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_197_io_data_1_in_valid = PENetwork_28_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_197_io_data_1_in_bits = PENetwork_28_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_197_io_data_0_in_valid = PENetwork_12_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_197_io_data_0_in_bits = PENetwork_12_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_197_io_sig_stat2trans = _T_1982_3; // @[pearray.scala 184:38]
  assign PE_198_clock = clock;
  assign PE_198_reset = reset;
  assign PE_198_io_data_2_in_valid = PENetwork_38_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_198_io_data_2_in_bits = PENetwork_38_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_198_io_data_1_in_valid = PENetwork_28_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_198_io_data_1_in_bits = PENetwork_28_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_198_io_data_0_in_valid = PENetwork_12_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_198_io_data_0_in_bits = PENetwork_12_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_198_io_sig_stat2trans = _T_1992_3; // @[pearray.scala 184:38]
  assign PE_199_clock = clock;
  assign PE_199_reset = reset;
  assign PE_199_io_data_2_in_valid = PENetwork_39_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_199_io_data_2_in_bits = PENetwork_39_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_199_io_data_1_in_valid = PENetwork_28_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_199_io_data_1_in_bits = PENetwork_28_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_199_io_data_0_in_valid = PENetwork_12_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_199_io_data_0_in_bits = PENetwork_12_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_199_io_sig_stat2trans = _T_2002_3; // @[pearray.scala 184:38]
  assign PE_200_clock = clock;
  assign PE_200_reset = reset;
  assign PE_200_io_data_2_in_valid = PENetwork_40_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_200_io_data_2_in_bits = PENetwork_40_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_200_io_data_1_in_valid = PENetwork_28_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_200_io_data_1_in_bits = PENetwork_28_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_200_io_data_0_in_valid = PENetwork_12_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_200_io_data_0_in_bits = PENetwork_12_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_200_io_sig_stat2trans = _T_2012_3; // @[pearray.scala 184:38]
  assign PE_201_clock = clock;
  assign PE_201_reset = reset;
  assign PE_201_io_data_2_in_valid = PENetwork_41_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_201_io_data_2_in_bits = PENetwork_41_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_201_io_data_1_in_valid = PENetwork_28_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_201_io_data_1_in_bits = PENetwork_28_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_201_io_data_0_in_valid = PENetwork_12_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_201_io_data_0_in_bits = PENetwork_12_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_201_io_sig_stat2trans = _T_2022_3; // @[pearray.scala 184:38]
  assign PE_202_clock = clock;
  assign PE_202_reset = reset;
  assign PE_202_io_data_2_in_valid = PENetwork_42_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_202_io_data_2_in_bits = PENetwork_42_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_202_io_data_1_in_valid = PENetwork_28_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_202_io_data_1_in_bits = PENetwork_28_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_202_io_data_0_in_valid = PENetwork_12_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_202_io_data_0_in_bits = PENetwork_12_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_202_io_sig_stat2trans = _T_2032_3; // @[pearray.scala 184:38]
  assign PE_203_clock = clock;
  assign PE_203_reset = reset;
  assign PE_203_io_data_2_in_valid = PENetwork_43_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_203_io_data_2_in_bits = PENetwork_43_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_203_io_data_1_in_valid = PENetwork_28_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_203_io_data_1_in_bits = PENetwork_28_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_203_io_data_0_in_valid = PENetwork_12_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_203_io_data_0_in_bits = PENetwork_12_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_203_io_sig_stat2trans = _T_2042_3; // @[pearray.scala 184:38]
  assign PE_204_clock = clock;
  assign PE_204_reset = reset;
  assign PE_204_io_data_2_in_valid = PENetwork_44_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_204_io_data_2_in_bits = PENetwork_44_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_204_io_data_1_in_valid = PENetwork_28_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_204_io_data_1_in_bits = PENetwork_28_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_204_io_data_0_in_valid = PENetwork_12_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_204_io_data_0_in_bits = PENetwork_12_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_204_io_sig_stat2trans = _T_2052_3; // @[pearray.scala 184:38]
  assign PE_205_clock = clock;
  assign PE_205_reset = reset;
  assign PE_205_io_data_2_in_valid = PENetwork_45_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_205_io_data_2_in_bits = PENetwork_45_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_205_io_data_1_in_valid = PENetwork_28_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_205_io_data_1_in_bits = PENetwork_28_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_205_io_data_0_in_valid = PENetwork_12_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_205_io_data_0_in_bits = PENetwork_12_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_205_io_sig_stat2trans = _T_2062_3; // @[pearray.scala 184:38]
  assign PE_206_clock = clock;
  assign PE_206_reset = reset;
  assign PE_206_io_data_2_in_valid = PENetwork_46_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_206_io_data_2_in_bits = PENetwork_46_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_206_io_data_1_in_valid = PENetwork_28_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_206_io_data_1_in_bits = PENetwork_28_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_206_io_data_0_in_valid = PENetwork_12_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_206_io_data_0_in_bits = PENetwork_12_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_206_io_sig_stat2trans = _T_2072_3; // @[pearray.scala 184:38]
  assign PE_207_clock = clock;
  assign PE_207_reset = reset;
  assign PE_207_io_data_2_in_valid = PENetwork_47_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_207_io_data_2_in_bits = PENetwork_47_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_207_io_data_1_in_valid = PENetwork_28_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_207_io_data_1_in_bits = PENetwork_28_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_207_io_data_0_in_valid = PENetwork_12_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_207_io_data_0_in_bits = PENetwork_12_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_207_io_sig_stat2trans = _T_2082_3; // @[pearray.scala 184:38]
  assign PE_208_clock = clock;
  assign PE_208_reset = reset;
  assign PE_208_io_data_2_in_valid = PENetwork_32_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_208_io_data_2_in_bits = PENetwork_32_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_208_io_data_1_in_valid = PENetwork_29_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_208_io_data_1_in_bits = PENetwork_29_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_208_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_208_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_208_io_sig_stat2trans = _T_2092_3; // @[pearray.scala 184:38]
  assign PE_209_clock = clock;
  assign PE_209_reset = reset;
  assign PE_209_io_data_2_in_valid = PENetwork_33_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_209_io_data_2_in_bits = PENetwork_33_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_209_io_data_1_in_valid = PENetwork_29_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_209_io_data_1_in_bits = PENetwork_29_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_209_io_data_0_in_valid = PENetwork_13_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_209_io_data_0_in_bits = PENetwork_13_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_209_io_sig_stat2trans = _T_2102_3; // @[pearray.scala 184:38]
  assign PE_210_clock = clock;
  assign PE_210_reset = reset;
  assign PE_210_io_data_2_in_valid = PENetwork_34_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_210_io_data_2_in_bits = PENetwork_34_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_210_io_data_1_in_valid = PENetwork_29_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_210_io_data_1_in_bits = PENetwork_29_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_210_io_data_0_in_valid = PENetwork_13_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_210_io_data_0_in_bits = PENetwork_13_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_210_io_sig_stat2trans = _T_2112_3; // @[pearray.scala 184:38]
  assign PE_211_clock = clock;
  assign PE_211_reset = reset;
  assign PE_211_io_data_2_in_valid = PENetwork_35_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_211_io_data_2_in_bits = PENetwork_35_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_211_io_data_1_in_valid = PENetwork_29_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_211_io_data_1_in_bits = PENetwork_29_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_211_io_data_0_in_valid = PENetwork_13_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_211_io_data_0_in_bits = PENetwork_13_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_211_io_sig_stat2trans = _T_2122_3; // @[pearray.scala 184:38]
  assign PE_212_clock = clock;
  assign PE_212_reset = reset;
  assign PE_212_io_data_2_in_valid = PENetwork_36_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_212_io_data_2_in_bits = PENetwork_36_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_212_io_data_1_in_valid = PENetwork_29_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_212_io_data_1_in_bits = PENetwork_29_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_212_io_data_0_in_valid = PENetwork_13_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_212_io_data_0_in_bits = PENetwork_13_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_212_io_sig_stat2trans = _T_2132_3; // @[pearray.scala 184:38]
  assign PE_213_clock = clock;
  assign PE_213_reset = reset;
  assign PE_213_io_data_2_in_valid = PENetwork_37_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_213_io_data_2_in_bits = PENetwork_37_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_213_io_data_1_in_valid = PENetwork_29_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_213_io_data_1_in_bits = PENetwork_29_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_213_io_data_0_in_valid = PENetwork_13_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_213_io_data_0_in_bits = PENetwork_13_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_213_io_sig_stat2trans = _T_2142_3; // @[pearray.scala 184:38]
  assign PE_214_clock = clock;
  assign PE_214_reset = reset;
  assign PE_214_io_data_2_in_valid = PENetwork_38_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_214_io_data_2_in_bits = PENetwork_38_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_214_io_data_1_in_valid = PENetwork_29_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_214_io_data_1_in_bits = PENetwork_29_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_214_io_data_0_in_valid = PENetwork_13_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_214_io_data_0_in_bits = PENetwork_13_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_214_io_sig_stat2trans = _T_2152_3; // @[pearray.scala 184:38]
  assign PE_215_clock = clock;
  assign PE_215_reset = reset;
  assign PE_215_io_data_2_in_valid = PENetwork_39_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_215_io_data_2_in_bits = PENetwork_39_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_215_io_data_1_in_valid = PENetwork_29_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_215_io_data_1_in_bits = PENetwork_29_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_215_io_data_0_in_valid = PENetwork_13_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_215_io_data_0_in_bits = PENetwork_13_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_215_io_sig_stat2trans = _T_2162_3; // @[pearray.scala 184:38]
  assign PE_216_clock = clock;
  assign PE_216_reset = reset;
  assign PE_216_io_data_2_in_valid = PENetwork_40_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_216_io_data_2_in_bits = PENetwork_40_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_216_io_data_1_in_valid = PENetwork_29_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_216_io_data_1_in_bits = PENetwork_29_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_216_io_data_0_in_valid = PENetwork_13_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_216_io_data_0_in_bits = PENetwork_13_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_216_io_sig_stat2trans = _T_2172_3; // @[pearray.scala 184:38]
  assign PE_217_clock = clock;
  assign PE_217_reset = reset;
  assign PE_217_io_data_2_in_valid = PENetwork_41_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_217_io_data_2_in_bits = PENetwork_41_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_217_io_data_1_in_valid = PENetwork_29_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_217_io_data_1_in_bits = PENetwork_29_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_217_io_data_0_in_valid = PENetwork_13_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_217_io_data_0_in_bits = PENetwork_13_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_217_io_sig_stat2trans = _T_2182_3; // @[pearray.scala 184:38]
  assign PE_218_clock = clock;
  assign PE_218_reset = reset;
  assign PE_218_io_data_2_in_valid = PENetwork_42_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_218_io_data_2_in_bits = PENetwork_42_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_218_io_data_1_in_valid = PENetwork_29_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_218_io_data_1_in_bits = PENetwork_29_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_218_io_data_0_in_valid = PENetwork_13_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_218_io_data_0_in_bits = PENetwork_13_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_218_io_sig_stat2trans = _T_2192_3; // @[pearray.scala 184:38]
  assign PE_219_clock = clock;
  assign PE_219_reset = reset;
  assign PE_219_io_data_2_in_valid = PENetwork_43_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_219_io_data_2_in_bits = PENetwork_43_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_219_io_data_1_in_valid = PENetwork_29_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_219_io_data_1_in_bits = PENetwork_29_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_219_io_data_0_in_valid = PENetwork_13_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_219_io_data_0_in_bits = PENetwork_13_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_219_io_sig_stat2trans = _T_2202_3; // @[pearray.scala 184:38]
  assign PE_220_clock = clock;
  assign PE_220_reset = reset;
  assign PE_220_io_data_2_in_valid = PENetwork_44_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_220_io_data_2_in_bits = PENetwork_44_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_220_io_data_1_in_valid = PENetwork_29_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_220_io_data_1_in_bits = PENetwork_29_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_220_io_data_0_in_valid = PENetwork_13_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_220_io_data_0_in_bits = PENetwork_13_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_220_io_sig_stat2trans = _T_2212_3; // @[pearray.scala 184:38]
  assign PE_221_clock = clock;
  assign PE_221_reset = reset;
  assign PE_221_io_data_2_in_valid = PENetwork_45_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_221_io_data_2_in_bits = PENetwork_45_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_221_io_data_1_in_valid = PENetwork_29_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_221_io_data_1_in_bits = PENetwork_29_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_221_io_data_0_in_valid = PENetwork_13_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_221_io_data_0_in_bits = PENetwork_13_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_221_io_sig_stat2trans = _T_2222_3; // @[pearray.scala 184:38]
  assign PE_222_clock = clock;
  assign PE_222_reset = reset;
  assign PE_222_io_data_2_in_valid = PENetwork_46_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_222_io_data_2_in_bits = PENetwork_46_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_222_io_data_1_in_valid = PENetwork_29_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_222_io_data_1_in_bits = PENetwork_29_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_222_io_data_0_in_valid = PENetwork_13_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_222_io_data_0_in_bits = PENetwork_13_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_222_io_sig_stat2trans = _T_2232_3; // @[pearray.scala 184:38]
  assign PE_223_clock = clock;
  assign PE_223_reset = reset;
  assign PE_223_io_data_2_in_valid = PENetwork_47_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_223_io_data_2_in_bits = PENetwork_47_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_223_io_data_1_in_valid = PENetwork_29_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_223_io_data_1_in_bits = PENetwork_29_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_223_io_data_0_in_valid = PENetwork_13_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_223_io_data_0_in_bits = PENetwork_13_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_223_io_sig_stat2trans = _T_2242_3; // @[pearray.scala 184:38]
  assign PE_224_clock = clock;
  assign PE_224_reset = reset;
  assign PE_224_io_data_2_in_valid = PENetwork_32_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_224_io_data_2_in_bits = PENetwork_32_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_224_io_data_1_in_valid = PENetwork_30_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_224_io_data_1_in_bits = PENetwork_30_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_224_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_224_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_224_io_sig_stat2trans = _T_2252_3; // @[pearray.scala 184:38]
  assign PE_225_clock = clock;
  assign PE_225_reset = reset;
  assign PE_225_io_data_2_in_valid = PENetwork_33_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_225_io_data_2_in_bits = PENetwork_33_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_225_io_data_1_in_valid = PENetwork_30_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_225_io_data_1_in_bits = PENetwork_30_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_225_io_data_0_in_valid = PENetwork_14_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_225_io_data_0_in_bits = PENetwork_14_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_225_io_sig_stat2trans = _T_2262_3; // @[pearray.scala 184:38]
  assign PE_226_clock = clock;
  assign PE_226_reset = reset;
  assign PE_226_io_data_2_in_valid = PENetwork_34_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_226_io_data_2_in_bits = PENetwork_34_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_226_io_data_1_in_valid = PENetwork_30_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_226_io_data_1_in_bits = PENetwork_30_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_226_io_data_0_in_valid = PENetwork_14_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_226_io_data_0_in_bits = PENetwork_14_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_226_io_sig_stat2trans = _T_2272_3; // @[pearray.scala 184:38]
  assign PE_227_clock = clock;
  assign PE_227_reset = reset;
  assign PE_227_io_data_2_in_valid = PENetwork_35_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_227_io_data_2_in_bits = PENetwork_35_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_227_io_data_1_in_valid = PENetwork_30_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_227_io_data_1_in_bits = PENetwork_30_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_227_io_data_0_in_valid = PENetwork_14_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_227_io_data_0_in_bits = PENetwork_14_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_227_io_sig_stat2trans = _T_2282_3; // @[pearray.scala 184:38]
  assign PE_228_clock = clock;
  assign PE_228_reset = reset;
  assign PE_228_io_data_2_in_valid = PENetwork_36_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_228_io_data_2_in_bits = PENetwork_36_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_228_io_data_1_in_valid = PENetwork_30_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_228_io_data_1_in_bits = PENetwork_30_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_228_io_data_0_in_valid = PENetwork_14_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_228_io_data_0_in_bits = PENetwork_14_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_228_io_sig_stat2trans = _T_2292_3; // @[pearray.scala 184:38]
  assign PE_229_clock = clock;
  assign PE_229_reset = reset;
  assign PE_229_io_data_2_in_valid = PENetwork_37_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_229_io_data_2_in_bits = PENetwork_37_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_229_io_data_1_in_valid = PENetwork_30_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_229_io_data_1_in_bits = PENetwork_30_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_229_io_data_0_in_valid = PENetwork_14_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_229_io_data_0_in_bits = PENetwork_14_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_229_io_sig_stat2trans = _T_2302_3; // @[pearray.scala 184:38]
  assign PE_230_clock = clock;
  assign PE_230_reset = reset;
  assign PE_230_io_data_2_in_valid = PENetwork_38_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_230_io_data_2_in_bits = PENetwork_38_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_230_io_data_1_in_valid = PENetwork_30_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_230_io_data_1_in_bits = PENetwork_30_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_230_io_data_0_in_valid = PENetwork_14_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_230_io_data_0_in_bits = PENetwork_14_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_230_io_sig_stat2trans = _T_2312_3; // @[pearray.scala 184:38]
  assign PE_231_clock = clock;
  assign PE_231_reset = reset;
  assign PE_231_io_data_2_in_valid = PENetwork_39_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_231_io_data_2_in_bits = PENetwork_39_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_231_io_data_1_in_valid = PENetwork_30_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_231_io_data_1_in_bits = PENetwork_30_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_231_io_data_0_in_valid = PENetwork_14_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_231_io_data_0_in_bits = PENetwork_14_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_231_io_sig_stat2trans = _T_2322_3; // @[pearray.scala 184:38]
  assign PE_232_clock = clock;
  assign PE_232_reset = reset;
  assign PE_232_io_data_2_in_valid = PENetwork_40_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_232_io_data_2_in_bits = PENetwork_40_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_232_io_data_1_in_valid = PENetwork_30_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_232_io_data_1_in_bits = PENetwork_30_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_232_io_data_0_in_valid = PENetwork_14_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_232_io_data_0_in_bits = PENetwork_14_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_232_io_sig_stat2trans = _T_2332_3; // @[pearray.scala 184:38]
  assign PE_233_clock = clock;
  assign PE_233_reset = reset;
  assign PE_233_io_data_2_in_valid = PENetwork_41_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_233_io_data_2_in_bits = PENetwork_41_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_233_io_data_1_in_valid = PENetwork_30_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_233_io_data_1_in_bits = PENetwork_30_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_233_io_data_0_in_valid = PENetwork_14_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_233_io_data_0_in_bits = PENetwork_14_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_233_io_sig_stat2trans = _T_2342_3; // @[pearray.scala 184:38]
  assign PE_234_clock = clock;
  assign PE_234_reset = reset;
  assign PE_234_io_data_2_in_valid = PENetwork_42_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_234_io_data_2_in_bits = PENetwork_42_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_234_io_data_1_in_valid = PENetwork_30_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_234_io_data_1_in_bits = PENetwork_30_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_234_io_data_0_in_valid = PENetwork_14_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_234_io_data_0_in_bits = PENetwork_14_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_234_io_sig_stat2trans = _T_2352_3; // @[pearray.scala 184:38]
  assign PE_235_clock = clock;
  assign PE_235_reset = reset;
  assign PE_235_io_data_2_in_valid = PENetwork_43_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_235_io_data_2_in_bits = PENetwork_43_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_235_io_data_1_in_valid = PENetwork_30_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_235_io_data_1_in_bits = PENetwork_30_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_235_io_data_0_in_valid = PENetwork_14_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_235_io_data_0_in_bits = PENetwork_14_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_235_io_sig_stat2trans = _T_2362_3; // @[pearray.scala 184:38]
  assign PE_236_clock = clock;
  assign PE_236_reset = reset;
  assign PE_236_io_data_2_in_valid = PENetwork_44_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_236_io_data_2_in_bits = PENetwork_44_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_236_io_data_1_in_valid = PENetwork_30_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_236_io_data_1_in_bits = PENetwork_30_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_236_io_data_0_in_valid = PENetwork_14_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_236_io_data_0_in_bits = PENetwork_14_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_236_io_sig_stat2trans = _T_2372_3; // @[pearray.scala 184:38]
  assign PE_237_clock = clock;
  assign PE_237_reset = reset;
  assign PE_237_io_data_2_in_valid = PENetwork_45_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_237_io_data_2_in_bits = PENetwork_45_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_237_io_data_1_in_valid = PENetwork_30_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_237_io_data_1_in_bits = PENetwork_30_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_237_io_data_0_in_valid = PENetwork_14_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_237_io_data_0_in_bits = PENetwork_14_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_237_io_sig_stat2trans = _T_2382_3; // @[pearray.scala 184:38]
  assign PE_238_clock = clock;
  assign PE_238_reset = reset;
  assign PE_238_io_data_2_in_valid = PENetwork_46_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_238_io_data_2_in_bits = PENetwork_46_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_238_io_data_1_in_valid = PENetwork_30_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_238_io_data_1_in_bits = PENetwork_30_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_238_io_data_0_in_valid = PENetwork_14_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_238_io_data_0_in_bits = PENetwork_14_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_238_io_sig_stat2trans = _T_2392_3; // @[pearray.scala 184:38]
  assign PE_239_clock = clock;
  assign PE_239_reset = reset;
  assign PE_239_io_data_2_in_valid = PENetwork_47_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_239_io_data_2_in_bits = PENetwork_47_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_239_io_data_1_in_valid = PENetwork_30_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_239_io_data_1_in_bits = PENetwork_30_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_239_io_data_0_in_valid = PENetwork_14_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_239_io_data_0_in_bits = PENetwork_14_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_239_io_sig_stat2trans = _T_2402_3; // @[pearray.scala 184:38]
  assign PE_240_clock = clock;
  assign PE_240_reset = reset;
  assign PE_240_io_data_2_in_valid = PENetwork_32_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_240_io_data_2_in_bits = PENetwork_32_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_240_io_data_1_in_valid = PENetwork_31_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_240_io_data_1_in_bits = PENetwork_31_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_240_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_240_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_240_io_sig_stat2trans = _T_2412_3; // @[pearray.scala 184:38]
  assign PE_241_clock = clock;
  assign PE_241_reset = reset;
  assign PE_241_io_data_2_in_valid = PENetwork_33_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_241_io_data_2_in_bits = PENetwork_33_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_241_io_data_1_in_valid = PENetwork_31_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_241_io_data_1_in_bits = PENetwork_31_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_241_io_data_0_in_valid = PENetwork_15_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_241_io_data_0_in_bits = PENetwork_15_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_241_io_sig_stat2trans = _T_2422_3; // @[pearray.scala 184:38]
  assign PE_242_clock = clock;
  assign PE_242_reset = reset;
  assign PE_242_io_data_2_in_valid = PENetwork_34_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_242_io_data_2_in_bits = PENetwork_34_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_242_io_data_1_in_valid = PENetwork_31_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_242_io_data_1_in_bits = PENetwork_31_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_242_io_data_0_in_valid = PENetwork_15_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_242_io_data_0_in_bits = PENetwork_15_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_242_io_sig_stat2trans = _T_2432_3; // @[pearray.scala 184:38]
  assign PE_243_clock = clock;
  assign PE_243_reset = reset;
  assign PE_243_io_data_2_in_valid = PENetwork_35_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_243_io_data_2_in_bits = PENetwork_35_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_243_io_data_1_in_valid = PENetwork_31_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_243_io_data_1_in_bits = PENetwork_31_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_243_io_data_0_in_valid = PENetwork_15_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_243_io_data_0_in_bits = PENetwork_15_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_243_io_sig_stat2trans = _T_2442_3; // @[pearray.scala 184:38]
  assign PE_244_clock = clock;
  assign PE_244_reset = reset;
  assign PE_244_io_data_2_in_valid = PENetwork_36_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_244_io_data_2_in_bits = PENetwork_36_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_244_io_data_1_in_valid = PENetwork_31_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_244_io_data_1_in_bits = PENetwork_31_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_244_io_data_0_in_valid = PENetwork_15_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_244_io_data_0_in_bits = PENetwork_15_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_244_io_sig_stat2trans = _T_2452_3; // @[pearray.scala 184:38]
  assign PE_245_clock = clock;
  assign PE_245_reset = reset;
  assign PE_245_io_data_2_in_valid = PENetwork_37_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_245_io_data_2_in_bits = PENetwork_37_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_245_io_data_1_in_valid = PENetwork_31_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_245_io_data_1_in_bits = PENetwork_31_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_245_io_data_0_in_valid = PENetwork_15_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_245_io_data_0_in_bits = PENetwork_15_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_245_io_sig_stat2trans = _T_2462_3; // @[pearray.scala 184:38]
  assign PE_246_clock = clock;
  assign PE_246_reset = reset;
  assign PE_246_io_data_2_in_valid = PENetwork_38_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_246_io_data_2_in_bits = PENetwork_38_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_246_io_data_1_in_valid = PENetwork_31_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_246_io_data_1_in_bits = PENetwork_31_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_246_io_data_0_in_valid = PENetwork_15_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_246_io_data_0_in_bits = PENetwork_15_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_246_io_sig_stat2trans = _T_2472_3; // @[pearray.scala 184:38]
  assign PE_247_clock = clock;
  assign PE_247_reset = reset;
  assign PE_247_io_data_2_in_valid = PENetwork_39_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_247_io_data_2_in_bits = PENetwork_39_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_247_io_data_1_in_valid = PENetwork_31_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_247_io_data_1_in_bits = PENetwork_31_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_247_io_data_0_in_valid = PENetwork_15_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_247_io_data_0_in_bits = PENetwork_15_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_247_io_sig_stat2trans = _T_2482_3; // @[pearray.scala 184:38]
  assign PE_248_clock = clock;
  assign PE_248_reset = reset;
  assign PE_248_io_data_2_in_valid = PENetwork_40_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_248_io_data_2_in_bits = PENetwork_40_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_248_io_data_1_in_valid = PENetwork_31_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_248_io_data_1_in_bits = PENetwork_31_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_248_io_data_0_in_valid = PENetwork_15_io_to_pes_8_in_valid; // @[pearray.scala 160:34]
  assign PE_248_io_data_0_in_bits = PENetwork_15_io_to_pes_8_in_bits; // @[pearray.scala 160:34]
  assign PE_248_io_sig_stat2trans = _T_2492_3; // @[pearray.scala 184:38]
  assign PE_249_clock = clock;
  assign PE_249_reset = reset;
  assign PE_249_io_data_2_in_valid = PENetwork_41_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_249_io_data_2_in_bits = PENetwork_41_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_249_io_data_1_in_valid = PENetwork_31_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_249_io_data_1_in_bits = PENetwork_31_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_249_io_data_0_in_valid = PENetwork_15_io_to_pes_9_in_valid; // @[pearray.scala 160:34]
  assign PE_249_io_data_0_in_bits = PENetwork_15_io_to_pes_9_in_bits; // @[pearray.scala 160:34]
  assign PE_249_io_sig_stat2trans = _T_2502_3; // @[pearray.scala 184:38]
  assign PE_250_clock = clock;
  assign PE_250_reset = reset;
  assign PE_250_io_data_2_in_valid = PENetwork_42_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_250_io_data_2_in_bits = PENetwork_42_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_250_io_data_1_in_valid = PENetwork_31_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_250_io_data_1_in_bits = PENetwork_31_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_250_io_data_0_in_valid = PENetwork_15_io_to_pes_10_in_valid; // @[pearray.scala 160:34]
  assign PE_250_io_data_0_in_bits = PENetwork_15_io_to_pes_10_in_bits; // @[pearray.scala 160:34]
  assign PE_250_io_sig_stat2trans = _T_2512_3; // @[pearray.scala 184:38]
  assign PE_251_clock = clock;
  assign PE_251_reset = reset;
  assign PE_251_io_data_2_in_valid = PENetwork_43_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_251_io_data_2_in_bits = PENetwork_43_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_251_io_data_1_in_valid = PENetwork_31_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_251_io_data_1_in_bits = PENetwork_31_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_251_io_data_0_in_valid = PENetwork_15_io_to_pes_11_in_valid; // @[pearray.scala 160:34]
  assign PE_251_io_data_0_in_bits = PENetwork_15_io_to_pes_11_in_bits; // @[pearray.scala 160:34]
  assign PE_251_io_sig_stat2trans = _T_2522_3; // @[pearray.scala 184:38]
  assign PE_252_clock = clock;
  assign PE_252_reset = reset;
  assign PE_252_io_data_2_in_valid = PENetwork_44_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_252_io_data_2_in_bits = PENetwork_44_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_252_io_data_1_in_valid = PENetwork_31_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_252_io_data_1_in_bits = PENetwork_31_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_252_io_data_0_in_valid = PENetwork_15_io_to_pes_12_in_valid; // @[pearray.scala 160:34]
  assign PE_252_io_data_0_in_bits = PENetwork_15_io_to_pes_12_in_bits; // @[pearray.scala 160:34]
  assign PE_252_io_sig_stat2trans = _T_2532_3; // @[pearray.scala 184:38]
  assign PE_253_clock = clock;
  assign PE_253_reset = reset;
  assign PE_253_io_data_2_in_valid = PENetwork_45_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_253_io_data_2_in_bits = PENetwork_45_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_253_io_data_1_in_valid = PENetwork_31_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_253_io_data_1_in_bits = PENetwork_31_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_253_io_data_0_in_valid = PENetwork_15_io_to_pes_13_in_valid; // @[pearray.scala 160:34]
  assign PE_253_io_data_0_in_bits = PENetwork_15_io_to_pes_13_in_bits; // @[pearray.scala 160:34]
  assign PE_253_io_sig_stat2trans = _T_2542_3; // @[pearray.scala 184:38]
  assign PE_254_clock = clock;
  assign PE_254_reset = reset;
  assign PE_254_io_data_2_in_valid = PENetwork_46_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_254_io_data_2_in_bits = PENetwork_46_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_254_io_data_1_in_valid = PENetwork_31_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_254_io_data_1_in_bits = PENetwork_31_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_254_io_data_0_in_valid = PENetwork_15_io_to_pes_14_in_valid; // @[pearray.scala 160:34]
  assign PE_254_io_data_0_in_bits = PENetwork_15_io_to_pes_14_in_bits; // @[pearray.scala 160:34]
  assign PE_254_io_sig_stat2trans = _T_2552_3; // @[pearray.scala 184:38]
  assign PE_255_clock = clock;
  assign PE_255_reset = reset;
  assign PE_255_io_data_2_in_valid = PENetwork_47_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_255_io_data_2_in_bits = PENetwork_47_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_255_io_data_1_in_valid = PENetwork_31_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_255_io_data_1_in_bits = PENetwork_31_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_255_io_data_0_in_valid = PENetwork_15_io_to_pes_15_in_valid; // @[pearray.scala 160:34]
  assign PE_255_io_data_0_in_bits = PENetwork_15_io_to_pes_15_in_bits; // @[pearray.scala 160:34]
  assign PE_255_io_sig_stat2trans = _T_2562_3; // @[pearray.scala 184:38]
  assign PENetwork_io_to_pes_0_out_valid = PE_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_0_out_bits = PE_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_1_out_valid = PE_1_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_1_out_bits = PE_1_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_2_out_valid = PE_2_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_2_out_bits = PE_2_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_3_out_valid = PE_3_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_3_out_bits = PE_3_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_4_out_valid = PE_4_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_4_out_bits = PE_4_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_5_out_valid = PE_5_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_5_out_bits = PE_5_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_6_out_valid = PE_6_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_6_out_bits = PE_6_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_7_out_valid = PE_7_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_7_out_bits = PE_7_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_8_out_valid = PE_8_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_8_out_bits = PE_8_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_9_out_valid = PE_9_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_9_out_bits = PE_9_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_10_out_valid = PE_10_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_10_out_bits = PE_10_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_11_out_valid = PE_11_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_11_out_bits = PE_11_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_12_out_valid = PE_12_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_12_out_bits = PE_12_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_13_out_valid = PE_13_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_13_out_bits = PE_13_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_14_out_valid = PE_14_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_14_out_bits = PE_14_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_15_out_valid = PE_15_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_15_out_bits = PE_15_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_0_out_valid = PE_16_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_0_out_bits = PE_16_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_1_out_valid = PE_17_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_1_out_bits = PE_17_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_2_out_valid = PE_18_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_2_out_bits = PE_18_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_3_out_valid = PE_19_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_3_out_bits = PE_19_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_4_out_valid = PE_20_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_4_out_bits = PE_20_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_5_out_valid = PE_21_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_5_out_bits = PE_21_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_6_out_valid = PE_22_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_6_out_bits = PE_22_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_7_out_valid = PE_23_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_7_out_bits = PE_23_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_8_out_valid = PE_24_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_8_out_bits = PE_24_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_9_out_valid = PE_25_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_9_out_bits = PE_25_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_10_out_valid = PE_26_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_10_out_bits = PE_26_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_11_out_valid = PE_27_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_11_out_bits = PE_27_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_12_out_valid = PE_28_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_12_out_bits = PE_28_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_13_out_valid = PE_29_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_13_out_bits = PE_29_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_14_out_valid = PE_30_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_14_out_bits = PE_30_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_15_out_valid = PE_31_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_15_out_bits = PE_31_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_0_out_valid = PE_32_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_0_out_bits = PE_32_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_1_out_valid = PE_33_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_1_out_bits = PE_33_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_2_out_valid = PE_34_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_2_out_bits = PE_34_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_3_out_valid = PE_35_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_3_out_bits = PE_35_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_4_out_valid = PE_36_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_4_out_bits = PE_36_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_5_out_valid = PE_37_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_5_out_bits = PE_37_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_6_out_valid = PE_38_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_6_out_bits = PE_38_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_7_out_valid = PE_39_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_7_out_bits = PE_39_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_8_out_valid = PE_40_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_8_out_bits = PE_40_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_9_out_valid = PE_41_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_9_out_bits = PE_41_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_10_out_valid = PE_42_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_10_out_bits = PE_42_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_11_out_valid = PE_43_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_11_out_bits = PE_43_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_12_out_valid = PE_44_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_12_out_bits = PE_44_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_13_out_valid = PE_45_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_13_out_bits = PE_45_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_14_out_valid = PE_46_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_14_out_bits = PE_46_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_15_out_valid = PE_47_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_15_out_bits = PE_47_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_0_out_valid = PE_48_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_0_out_bits = PE_48_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_1_out_valid = PE_49_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_1_out_bits = PE_49_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_2_out_valid = PE_50_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_2_out_bits = PE_50_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_3_out_valid = PE_51_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_3_out_bits = PE_51_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_4_out_valid = PE_52_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_4_out_bits = PE_52_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_5_out_valid = PE_53_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_5_out_bits = PE_53_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_6_out_valid = PE_54_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_6_out_bits = PE_54_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_7_out_valid = PE_55_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_7_out_bits = PE_55_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_8_out_valid = PE_56_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_8_out_bits = PE_56_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_9_out_valid = PE_57_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_9_out_bits = PE_57_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_10_out_valid = PE_58_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_10_out_bits = PE_58_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_11_out_valid = PE_59_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_11_out_bits = PE_59_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_12_out_valid = PE_60_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_12_out_bits = PE_60_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_13_out_valid = PE_61_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_13_out_bits = PE_61_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_14_out_valid = PE_62_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_14_out_bits = PE_62_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_15_out_valid = PE_63_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_15_out_bits = PE_63_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_0_out_valid = PE_64_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_0_out_bits = PE_64_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_1_out_valid = PE_65_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_1_out_bits = PE_65_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_2_out_valid = PE_66_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_2_out_bits = PE_66_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_3_out_valid = PE_67_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_3_out_bits = PE_67_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_4_out_valid = PE_68_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_4_out_bits = PE_68_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_5_out_valid = PE_69_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_5_out_bits = PE_69_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_6_out_valid = PE_70_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_6_out_bits = PE_70_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_7_out_valid = PE_71_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_7_out_bits = PE_71_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_8_out_valid = PE_72_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_8_out_bits = PE_72_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_9_out_valid = PE_73_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_9_out_bits = PE_73_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_10_out_valid = PE_74_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_10_out_bits = PE_74_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_11_out_valid = PE_75_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_11_out_bits = PE_75_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_12_out_valid = PE_76_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_12_out_bits = PE_76_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_13_out_valid = PE_77_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_13_out_bits = PE_77_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_14_out_valid = PE_78_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_14_out_bits = PE_78_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_15_out_valid = PE_79_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_15_out_bits = PE_79_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_0_out_valid = PE_80_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_0_out_bits = PE_80_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_1_out_valid = PE_81_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_1_out_bits = PE_81_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_2_out_valid = PE_82_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_2_out_bits = PE_82_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_3_out_valid = PE_83_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_3_out_bits = PE_83_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_4_out_valid = PE_84_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_4_out_bits = PE_84_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_5_out_valid = PE_85_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_5_out_bits = PE_85_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_6_out_valid = PE_86_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_6_out_bits = PE_86_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_7_out_valid = PE_87_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_7_out_bits = PE_87_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_8_out_valid = PE_88_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_8_out_bits = PE_88_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_9_out_valid = PE_89_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_9_out_bits = PE_89_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_10_out_valid = PE_90_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_10_out_bits = PE_90_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_11_out_valid = PE_91_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_11_out_bits = PE_91_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_12_out_valid = PE_92_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_12_out_bits = PE_92_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_13_out_valid = PE_93_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_13_out_bits = PE_93_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_14_out_valid = PE_94_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_14_out_bits = PE_94_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_15_out_valid = PE_95_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_15_out_bits = PE_95_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_0_out_valid = PE_96_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_0_out_bits = PE_96_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_1_out_valid = PE_97_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_1_out_bits = PE_97_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_2_out_valid = PE_98_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_2_out_bits = PE_98_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_3_out_valid = PE_99_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_3_out_bits = PE_99_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_4_out_valid = PE_100_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_4_out_bits = PE_100_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_5_out_valid = PE_101_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_5_out_bits = PE_101_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_6_out_valid = PE_102_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_6_out_bits = PE_102_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_7_out_valid = PE_103_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_7_out_bits = PE_103_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_8_out_valid = PE_104_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_8_out_bits = PE_104_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_9_out_valid = PE_105_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_9_out_bits = PE_105_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_10_out_valid = PE_106_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_10_out_bits = PE_106_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_11_out_valid = PE_107_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_11_out_bits = PE_107_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_12_out_valid = PE_108_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_12_out_bits = PE_108_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_13_out_valid = PE_109_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_13_out_bits = PE_109_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_14_out_valid = PE_110_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_14_out_bits = PE_110_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_15_out_valid = PE_111_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_15_out_bits = PE_111_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_0_out_valid = PE_112_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_0_out_bits = PE_112_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_1_out_valid = PE_113_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_1_out_bits = PE_113_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_2_out_valid = PE_114_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_2_out_bits = PE_114_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_3_out_valid = PE_115_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_3_out_bits = PE_115_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_4_out_valid = PE_116_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_4_out_bits = PE_116_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_5_out_valid = PE_117_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_5_out_bits = PE_117_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_6_out_valid = PE_118_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_6_out_bits = PE_118_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_7_out_valid = PE_119_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_7_out_bits = PE_119_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_8_out_valid = PE_120_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_8_out_bits = PE_120_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_9_out_valid = PE_121_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_9_out_bits = PE_121_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_10_out_valid = PE_122_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_10_out_bits = PE_122_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_11_out_valid = PE_123_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_11_out_bits = PE_123_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_12_out_valid = PE_124_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_12_out_bits = PE_124_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_13_out_valid = PE_125_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_13_out_bits = PE_125_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_14_out_valid = PE_126_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_14_out_bits = PE_126_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_15_out_valid = PE_127_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_15_out_bits = PE_127_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_0_out_valid = PE_128_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_0_out_bits = PE_128_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_1_out_valid = PE_129_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_1_out_bits = PE_129_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_2_out_valid = PE_130_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_2_out_bits = PE_130_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_3_out_valid = PE_131_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_3_out_bits = PE_131_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_4_out_valid = PE_132_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_4_out_bits = PE_132_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_5_out_valid = PE_133_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_5_out_bits = PE_133_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_6_out_valid = PE_134_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_6_out_bits = PE_134_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_7_out_valid = PE_135_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_7_out_bits = PE_135_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_8_out_valid = PE_136_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_8_out_bits = PE_136_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_9_out_valid = PE_137_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_9_out_bits = PE_137_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_10_out_valid = PE_138_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_10_out_bits = PE_138_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_11_out_valid = PE_139_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_11_out_bits = PE_139_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_12_out_valid = PE_140_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_12_out_bits = PE_140_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_13_out_valid = PE_141_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_13_out_bits = PE_141_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_14_out_valid = PE_142_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_14_out_bits = PE_142_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_15_out_valid = PE_143_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_15_out_bits = PE_143_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_0_out_valid = PE_144_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_0_out_bits = PE_144_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_1_out_valid = PE_145_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_1_out_bits = PE_145_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_2_out_valid = PE_146_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_2_out_bits = PE_146_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_3_out_valid = PE_147_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_3_out_bits = PE_147_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_4_out_valid = PE_148_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_4_out_bits = PE_148_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_5_out_valid = PE_149_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_5_out_bits = PE_149_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_6_out_valid = PE_150_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_6_out_bits = PE_150_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_7_out_valid = PE_151_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_7_out_bits = PE_151_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_8_out_valid = PE_152_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_8_out_bits = PE_152_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_9_out_valid = PE_153_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_9_out_bits = PE_153_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_10_out_valid = PE_154_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_10_out_bits = PE_154_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_11_out_valid = PE_155_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_11_out_bits = PE_155_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_12_out_valid = PE_156_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_12_out_bits = PE_156_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_13_out_valid = PE_157_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_13_out_bits = PE_157_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_14_out_valid = PE_158_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_14_out_bits = PE_158_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_15_out_valid = PE_159_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_15_out_bits = PE_159_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_0_out_valid = PE_160_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_0_out_bits = PE_160_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_1_out_valid = PE_161_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_1_out_bits = PE_161_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_2_out_valid = PE_162_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_2_out_bits = PE_162_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_3_out_valid = PE_163_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_3_out_bits = PE_163_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_4_out_valid = PE_164_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_4_out_bits = PE_164_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_5_out_valid = PE_165_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_5_out_bits = PE_165_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_6_out_valid = PE_166_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_6_out_bits = PE_166_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_7_out_valid = PE_167_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_7_out_bits = PE_167_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_8_out_valid = PE_168_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_8_out_bits = PE_168_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_9_out_valid = PE_169_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_9_out_bits = PE_169_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_10_out_valid = PE_170_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_10_out_bits = PE_170_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_11_out_valid = PE_171_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_11_out_bits = PE_171_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_12_out_valid = PE_172_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_12_out_bits = PE_172_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_13_out_valid = PE_173_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_13_out_bits = PE_173_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_14_out_valid = PE_174_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_14_out_bits = PE_174_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_15_out_valid = PE_175_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_15_out_bits = PE_175_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_0_out_valid = PE_176_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_0_out_bits = PE_176_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_1_out_valid = PE_177_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_1_out_bits = PE_177_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_2_out_valid = PE_178_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_2_out_bits = PE_178_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_3_out_valid = PE_179_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_3_out_bits = PE_179_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_4_out_valid = PE_180_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_4_out_bits = PE_180_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_5_out_valid = PE_181_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_5_out_bits = PE_181_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_6_out_valid = PE_182_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_6_out_bits = PE_182_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_7_out_valid = PE_183_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_7_out_bits = PE_183_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_8_out_valid = PE_184_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_8_out_bits = PE_184_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_9_out_valid = PE_185_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_9_out_bits = PE_185_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_10_out_valid = PE_186_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_10_out_bits = PE_186_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_11_out_valid = PE_187_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_11_out_bits = PE_187_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_12_out_valid = PE_188_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_12_out_bits = PE_188_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_13_out_valid = PE_189_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_13_out_bits = PE_189_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_14_out_valid = PE_190_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_14_out_bits = PE_190_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_15_out_valid = PE_191_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_15_out_bits = PE_191_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_0_out_valid = PE_192_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_0_out_bits = PE_192_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_1_out_valid = PE_193_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_1_out_bits = PE_193_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_2_out_valid = PE_194_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_2_out_bits = PE_194_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_3_out_valid = PE_195_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_3_out_bits = PE_195_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_4_out_valid = PE_196_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_4_out_bits = PE_196_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_5_out_valid = PE_197_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_5_out_bits = PE_197_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_6_out_valid = PE_198_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_6_out_bits = PE_198_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_7_out_valid = PE_199_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_7_out_bits = PE_199_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_8_out_valid = PE_200_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_8_out_bits = PE_200_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_9_out_valid = PE_201_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_9_out_bits = PE_201_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_10_out_valid = PE_202_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_10_out_bits = PE_202_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_11_out_valid = PE_203_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_11_out_bits = PE_203_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_12_out_valid = PE_204_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_12_out_bits = PE_204_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_13_out_valid = PE_205_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_13_out_bits = PE_205_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_14_out_valid = PE_206_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_14_out_bits = PE_206_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_15_out_valid = PE_207_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_15_out_bits = PE_207_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_0_out_valid = PE_208_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_0_out_bits = PE_208_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_1_out_valid = PE_209_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_1_out_bits = PE_209_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_2_out_valid = PE_210_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_2_out_bits = PE_210_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_3_out_valid = PE_211_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_3_out_bits = PE_211_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_4_out_valid = PE_212_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_4_out_bits = PE_212_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_5_out_valid = PE_213_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_5_out_bits = PE_213_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_6_out_valid = PE_214_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_6_out_bits = PE_214_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_7_out_valid = PE_215_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_7_out_bits = PE_215_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_8_out_valid = PE_216_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_8_out_bits = PE_216_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_9_out_valid = PE_217_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_9_out_bits = PE_217_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_10_out_valid = PE_218_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_10_out_bits = PE_218_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_11_out_valid = PE_219_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_11_out_bits = PE_219_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_12_out_valid = PE_220_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_12_out_bits = PE_220_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_13_out_valid = PE_221_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_13_out_bits = PE_221_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_14_out_valid = PE_222_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_14_out_bits = PE_222_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_15_out_valid = PE_223_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_15_out_bits = PE_223_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_0_out_valid = PE_224_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_0_out_bits = PE_224_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_1_out_valid = PE_225_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_1_out_bits = PE_225_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_2_out_valid = PE_226_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_2_out_bits = PE_226_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_3_out_valid = PE_227_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_3_out_bits = PE_227_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_4_out_valid = PE_228_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_4_out_bits = PE_228_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_5_out_valid = PE_229_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_5_out_bits = PE_229_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_6_out_valid = PE_230_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_6_out_bits = PE_230_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_7_out_valid = PE_231_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_7_out_bits = PE_231_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_8_out_valid = PE_232_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_8_out_bits = PE_232_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_9_out_valid = PE_233_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_9_out_bits = PE_233_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_10_out_valid = PE_234_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_10_out_bits = PE_234_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_11_out_valid = PE_235_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_11_out_bits = PE_235_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_12_out_valid = PE_236_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_12_out_bits = PE_236_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_13_out_valid = PE_237_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_13_out_bits = PE_237_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_14_out_valid = PE_238_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_14_out_bits = PE_238_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_15_out_valid = PE_239_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_15_out_bits = PE_239_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_0_out_valid = PE_240_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_0_out_bits = PE_240_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_1_out_valid = PE_241_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_1_out_bits = PE_241_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_2_out_valid = PE_242_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_2_out_bits = PE_242_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_3_out_valid = PE_243_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_3_out_bits = PE_243_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_4_out_valid = PE_244_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_4_out_bits = PE_244_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_5_out_valid = PE_245_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_5_out_bits = PE_245_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_6_out_valid = PE_246_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_6_out_bits = PE_246_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_7_out_valid = PE_247_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_7_out_bits = PE_247_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_8_out_valid = PE_248_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_8_out_bits = PE_248_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_9_out_valid = PE_249_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_9_out_bits = PE_249_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_10_out_valid = PE_250_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_10_out_bits = PE_250_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_11_out_valid = PE_251_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_11_out_bits = PE_251_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_12_out_valid = PE_252_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_12_out_bits = PE_252_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_13_out_valid = PE_253_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_13_out_bits = PE_253_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_14_out_valid = PE_254_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_14_out_bits = PE_254_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_15_out_valid = PE_255_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_15_out_bits = PE_255_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_0_out_valid = PE_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_0_out_bits = PE_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_1_out_valid = PE_1_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_1_out_bits = PE_1_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_2_out_valid = PE_2_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_2_out_bits = PE_2_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_3_out_valid = PE_3_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_3_out_bits = PE_3_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_4_out_valid = PE_4_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_4_out_bits = PE_4_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_5_out_valid = PE_5_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_5_out_bits = PE_5_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_6_out_valid = PE_6_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_6_out_bits = PE_6_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_7_out_valid = PE_7_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_7_out_bits = PE_7_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_8_out_valid = PE_8_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_8_out_bits = PE_8_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_9_out_valid = PE_9_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_9_out_bits = PE_9_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_10_out_valid = PE_10_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_10_out_bits = PE_10_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_11_out_valid = PE_11_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_11_out_bits = PE_11_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_12_out_valid = PE_12_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_12_out_bits = PE_12_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_13_out_valid = PE_13_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_13_out_bits = PE_13_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_14_out_valid = PE_14_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_14_out_bits = PE_14_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_mem_valid = MemController_16_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_16_io_to_mem_bits = MemController_16_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_17_io_to_pes_0_out_valid = PE_16_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_0_out_bits = PE_16_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_1_out_valid = PE_17_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_1_out_bits = PE_17_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_2_out_valid = PE_18_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_2_out_bits = PE_18_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_3_out_valid = PE_19_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_3_out_bits = PE_19_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_4_out_valid = PE_20_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_4_out_bits = PE_20_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_5_out_valid = PE_21_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_5_out_bits = PE_21_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_6_out_valid = PE_22_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_6_out_bits = PE_22_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_7_out_valid = PE_23_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_7_out_bits = PE_23_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_8_out_valid = PE_24_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_8_out_bits = PE_24_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_9_out_valid = PE_25_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_9_out_bits = PE_25_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_10_out_valid = PE_26_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_10_out_bits = PE_26_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_11_out_valid = PE_27_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_11_out_bits = PE_27_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_12_out_valid = PE_28_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_12_out_bits = PE_28_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_13_out_valid = PE_29_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_13_out_bits = PE_29_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_14_out_valid = PE_30_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_14_out_bits = PE_30_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_mem_valid = MemController_17_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_17_io_to_mem_bits = MemController_17_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_18_io_to_pes_0_out_valid = PE_32_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_0_out_bits = PE_32_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_1_out_valid = PE_33_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_1_out_bits = PE_33_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_2_out_valid = PE_34_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_2_out_bits = PE_34_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_3_out_valid = PE_35_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_3_out_bits = PE_35_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_4_out_valid = PE_36_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_4_out_bits = PE_36_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_5_out_valid = PE_37_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_5_out_bits = PE_37_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_6_out_valid = PE_38_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_6_out_bits = PE_38_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_7_out_valid = PE_39_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_7_out_bits = PE_39_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_8_out_valid = PE_40_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_8_out_bits = PE_40_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_9_out_valid = PE_41_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_9_out_bits = PE_41_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_10_out_valid = PE_42_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_10_out_bits = PE_42_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_11_out_valid = PE_43_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_11_out_bits = PE_43_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_12_out_valid = PE_44_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_12_out_bits = PE_44_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_13_out_valid = PE_45_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_13_out_bits = PE_45_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_14_out_valid = PE_46_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_14_out_bits = PE_46_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_mem_valid = MemController_18_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_18_io_to_mem_bits = MemController_18_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_19_io_to_pes_0_out_valid = PE_48_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_0_out_bits = PE_48_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_1_out_valid = PE_49_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_1_out_bits = PE_49_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_2_out_valid = PE_50_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_2_out_bits = PE_50_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_3_out_valid = PE_51_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_3_out_bits = PE_51_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_4_out_valid = PE_52_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_4_out_bits = PE_52_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_5_out_valid = PE_53_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_5_out_bits = PE_53_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_6_out_valid = PE_54_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_6_out_bits = PE_54_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_7_out_valid = PE_55_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_7_out_bits = PE_55_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_8_out_valid = PE_56_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_8_out_bits = PE_56_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_9_out_valid = PE_57_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_9_out_bits = PE_57_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_10_out_valid = PE_58_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_10_out_bits = PE_58_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_11_out_valid = PE_59_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_11_out_bits = PE_59_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_12_out_valid = PE_60_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_12_out_bits = PE_60_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_13_out_valid = PE_61_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_13_out_bits = PE_61_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_14_out_valid = PE_62_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_14_out_bits = PE_62_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_mem_valid = MemController_19_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_19_io_to_mem_bits = MemController_19_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_20_io_to_pes_0_out_valid = PE_64_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_0_out_bits = PE_64_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_1_out_valid = PE_65_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_1_out_bits = PE_65_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_2_out_valid = PE_66_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_2_out_bits = PE_66_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_3_out_valid = PE_67_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_3_out_bits = PE_67_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_4_out_valid = PE_68_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_4_out_bits = PE_68_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_5_out_valid = PE_69_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_5_out_bits = PE_69_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_6_out_valid = PE_70_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_6_out_bits = PE_70_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_7_out_valid = PE_71_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_7_out_bits = PE_71_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_8_out_valid = PE_72_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_8_out_bits = PE_72_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_9_out_valid = PE_73_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_9_out_bits = PE_73_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_10_out_valid = PE_74_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_10_out_bits = PE_74_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_11_out_valid = PE_75_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_11_out_bits = PE_75_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_12_out_valid = PE_76_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_12_out_bits = PE_76_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_13_out_valid = PE_77_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_13_out_bits = PE_77_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_14_out_valid = PE_78_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_14_out_bits = PE_78_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_mem_valid = MemController_20_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_20_io_to_mem_bits = MemController_20_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_21_io_to_pes_0_out_valid = PE_80_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_0_out_bits = PE_80_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_1_out_valid = PE_81_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_1_out_bits = PE_81_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_2_out_valid = PE_82_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_2_out_bits = PE_82_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_3_out_valid = PE_83_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_3_out_bits = PE_83_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_4_out_valid = PE_84_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_4_out_bits = PE_84_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_5_out_valid = PE_85_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_5_out_bits = PE_85_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_6_out_valid = PE_86_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_6_out_bits = PE_86_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_7_out_valid = PE_87_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_7_out_bits = PE_87_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_8_out_valid = PE_88_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_8_out_bits = PE_88_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_9_out_valid = PE_89_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_9_out_bits = PE_89_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_10_out_valid = PE_90_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_10_out_bits = PE_90_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_11_out_valid = PE_91_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_11_out_bits = PE_91_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_12_out_valid = PE_92_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_12_out_bits = PE_92_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_13_out_valid = PE_93_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_13_out_bits = PE_93_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_14_out_valid = PE_94_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_14_out_bits = PE_94_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_mem_valid = MemController_21_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_21_io_to_mem_bits = MemController_21_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_22_io_to_pes_0_out_valid = PE_96_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_0_out_bits = PE_96_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_1_out_valid = PE_97_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_1_out_bits = PE_97_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_2_out_valid = PE_98_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_2_out_bits = PE_98_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_3_out_valid = PE_99_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_3_out_bits = PE_99_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_4_out_valid = PE_100_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_4_out_bits = PE_100_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_5_out_valid = PE_101_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_5_out_bits = PE_101_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_6_out_valid = PE_102_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_6_out_bits = PE_102_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_7_out_valid = PE_103_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_7_out_bits = PE_103_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_8_out_valid = PE_104_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_8_out_bits = PE_104_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_9_out_valid = PE_105_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_9_out_bits = PE_105_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_10_out_valid = PE_106_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_10_out_bits = PE_106_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_11_out_valid = PE_107_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_11_out_bits = PE_107_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_12_out_valid = PE_108_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_12_out_bits = PE_108_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_13_out_valid = PE_109_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_13_out_bits = PE_109_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_14_out_valid = PE_110_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_14_out_bits = PE_110_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_mem_valid = MemController_22_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_22_io_to_mem_bits = MemController_22_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_23_io_to_pes_0_out_valid = PE_112_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_0_out_bits = PE_112_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_1_out_valid = PE_113_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_1_out_bits = PE_113_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_2_out_valid = PE_114_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_2_out_bits = PE_114_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_3_out_valid = PE_115_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_3_out_bits = PE_115_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_4_out_valid = PE_116_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_4_out_bits = PE_116_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_5_out_valid = PE_117_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_5_out_bits = PE_117_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_6_out_valid = PE_118_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_6_out_bits = PE_118_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_7_out_valid = PE_119_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_7_out_bits = PE_119_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_8_out_valid = PE_120_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_8_out_bits = PE_120_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_9_out_valid = PE_121_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_9_out_bits = PE_121_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_10_out_valid = PE_122_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_10_out_bits = PE_122_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_11_out_valid = PE_123_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_11_out_bits = PE_123_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_12_out_valid = PE_124_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_12_out_bits = PE_124_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_13_out_valid = PE_125_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_13_out_bits = PE_125_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_14_out_valid = PE_126_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_14_out_bits = PE_126_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_mem_valid = MemController_23_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_23_io_to_mem_bits = MemController_23_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_24_io_to_pes_0_out_valid = PE_128_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_0_out_bits = PE_128_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_1_out_valid = PE_129_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_1_out_bits = PE_129_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_2_out_valid = PE_130_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_2_out_bits = PE_130_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_3_out_valid = PE_131_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_3_out_bits = PE_131_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_4_out_valid = PE_132_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_4_out_bits = PE_132_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_5_out_valid = PE_133_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_5_out_bits = PE_133_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_6_out_valid = PE_134_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_6_out_bits = PE_134_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_7_out_valid = PE_135_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_7_out_bits = PE_135_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_8_out_valid = PE_136_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_8_out_bits = PE_136_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_9_out_valid = PE_137_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_9_out_bits = PE_137_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_10_out_valid = PE_138_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_10_out_bits = PE_138_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_11_out_valid = PE_139_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_11_out_bits = PE_139_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_12_out_valid = PE_140_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_12_out_bits = PE_140_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_13_out_valid = PE_141_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_13_out_bits = PE_141_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_14_out_valid = PE_142_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_pes_14_out_bits = PE_142_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_24_io_to_mem_valid = MemController_24_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_24_io_to_mem_bits = MemController_24_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_25_io_to_pes_0_out_valid = PE_144_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_0_out_bits = PE_144_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_1_out_valid = PE_145_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_1_out_bits = PE_145_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_2_out_valid = PE_146_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_2_out_bits = PE_146_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_3_out_valid = PE_147_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_3_out_bits = PE_147_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_4_out_valid = PE_148_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_4_out_bits = PE_148_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_5_out_valid = PE_149_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_5_out_bits = PE_149_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_6_out_valid = PE_150_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_6_out_bits = PE_150_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_7_out_valid = PE_151_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_7_out_bits = PE_151_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_8_out_valid = PE_152_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_8_out_bits = PE_152_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_9_out_valid = PE_153_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_9_out_bits = PE_153_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_10_out_valid = PE_154_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_10_out_bits = PE_154_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_11_out_valid = PE_155_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_11_out_bits = PE_155_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_12_out_valid = PE_156_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_12_out_bits = PE_156_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_13_out_valid = PE_157_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_13_out_bits = PE_157_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_14_out_valid = PE_158_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_pes_14_out_bits = PE_158_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_25_io_to_mem_valid = MemController_25_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_25_io_to_mem_bits = MemController_25_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_26_io_to_pes_0_out_valid = PE_160_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_0_out_bits = PE_160_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_1_out_valid = PE_161_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_1_out_bits = PE_161_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_2_out_valid = PE_162_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_2_out_bits = PE_162_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_3_out_valid = PE_163_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_3_out_bits = PE_163_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_4_out_valid = PE_164_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_4_out_bits = PE_164_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_5_out_valid = PE_165_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_5_out_bits = PE_165_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_6_out_valid = PE_166_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_6_out_bits = PE_166_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_7_out_valid = PE_167_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_7_out_bits = PE_167_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_8_out_valid = PE_168_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_8_out_bits = PE_168_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_9_out_valid = PE_169_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_9_out_bits = PE_169_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_10_out_valid = PE_170_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_10_out_bits = PE_170_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_11_out_valid = PE_171_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_11_out_bits = PE_171_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_12_out_valid = PE_172_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_12_out_bits = PE_172_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_13_out_valid = PE_173_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_13_out_bits = PE_173_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_14_out_valid = PE_174_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_pes_14_out_bits = PE_174_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_26_io_to_mem_valid = MemController_26_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_26_io_to_mem_bits = MemController_26_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_27_io_to_pes_0_out_valid = PE_176_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_0_out_bits = PE_176_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_1_out_valid = PE_177_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_1_out_bits = PE_177_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_2_out_valid = PE_178_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_2_out_bits = PE_178_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_3_out_valid = PE_179_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_3_out_bits = PE_179_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_4_out_valid = PE_180_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_4_out_bits = PE_180_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_5_out_valid = PE_181_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_5_out_bits = PE_181_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_6_out_valid = PE_182_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_6_out_bits = PE_182_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_7_out_valid = PE_183_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_7_out_bits = PE_183_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_8_out_valid = PE_184_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_8_out_bits = PE_184_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_9_out_valid = PE_185_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_9_out_bits = PE_185_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_10_out_valid = PE_186_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_10_out_bits = PE_186_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_11_out_valid = PE_187_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_11_out_bits = PE_187_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_12_out_valid = PE_188_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_12_out_bits = PE_188_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_13_out_valid = PE_189_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_13_out_bits = PE_189_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_14_out_valid = PE_190_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_pes_14_out_bits = PE_190_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_27_io_to_mem_valid = MemController_27_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_27_io_to_mem_bits = MemController_27_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_28_io_to_pes_0_out_valid = PE_192_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_0_out_bits = PE_192_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_1_out_valid = PE_193_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_1_out_bits = PE_193_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_2_out_valid = PE_194_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_2_out_bits = PE_194_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_3_out_valid = PE_195_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_3_out_bits = PE_195_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_4_out_valid = PE_196_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_4_out_bits = PE_196_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_5_out_valid = PE_197_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_5_out_bits = PE_197_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_6_out_valid = PE_198_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_6_out_bits = PE_198_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_7_out_valid = PE_199_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_7_out_bits = PE_199_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_8_out_valid = PE_200_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_8_out_bits = PE_200_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_9_out_valid = PE_201_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_9_out_bits = PE_201_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_10_out_valid = PE_202_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_10_out_bits = PE_202_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_11_out_valid = PE_203_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_11_out_bits = PE_203_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_12_out_valid = PE_204_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_12_out_bits = PE_204_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_13_out_valid = PE_205_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_13_out_bits = PE_205_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_14_out_valid = PE_206_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_pes_14_out_bits = PE_206_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_28_io_to_mem_valid = MemController_28_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_28_io_to_mem_bits = MemController_28_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_29_io_to_pes_0_out_valid = PE_208_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_0_out_bits = PE_208_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_1_out_valid = PE_209_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_1_out_bits = PE_209_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_2_out_valid = PE_210_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_2_out_bits = PE_210_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_3_out_valid = PE_211_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_3_out_bits = PE_211_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_4_out_valid = PE_212_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_4_out_bits = PE_212_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_5_out_valid = PE_213_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_5_out_bits = PE_213_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_6_out_valid = PE_214_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_6_out_bits = PE_214_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_7_out_valid = PE_215_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_7_out_bits = PE_215_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_8_out_valid = PE_216_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_8_out_bits = PE_216_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_9_out_valid = PE_217_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_9_out_bits = PE_217_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_10_out_valid = PE_218_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_10_out_bits = PE_218_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_11_out_valid = PE_219_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_11_out_bits = PE_219_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_12_out_valid = PE_220_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_12_out_bits = PE_220_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_13_out_valid = PE_221_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_13_out_bits = PE_221_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_14_out_valid = PE_222_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_pes_14_out_bits = PE_222_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_29_io_to_mem_valid = MemController_29_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_29_io_to_mem_bits = MemController_29_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_30_io_to_pes_0_out_valid = PE_224_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_0_out_bits = PE_224_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_1_out_valid = PE_225_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_1_out_bits = PE_225_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_2_out_valid = PE_226_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_2_out_bits = PE_226_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_3_out_valid = PE_227_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_3_out_bits = PE_227_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_4_out_valid = PE_228_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_4_out_bits = PE_228_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_5_out_valid = PE_229_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_5_out_bits = PE_229_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_6_out_valid = PE_230_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_6_out_bits = PE_230_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_7_out_valid = PE_231_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_7_out_bits = PE_231_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_8_out_valid = PE_232_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_8_out_bits = PE_232_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_9_out_valid = PE_233_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_9_out_bits = PE_233_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_10_out_valid = PE_234_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_10_out_bits = PE_234_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_11_out_valid = PE_235_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_11_out_bits = PE_235_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_12_out_valid = PE_236_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_12_out_bits = PE_236_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_13_out_valid = PE_237_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_13_out_bits = PE_237_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_14_out_valid = PE_238_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_pes_14_out_bits = PE_238_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_30_io_to_mem_valid = MemController_30_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_30_io_to_mem_bits = MemController_30_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_31_io_to_pes_0_out_valid = PE_240_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_0_out_bits = PE_240_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_1_out_valid = PE_241_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_1_out_bits = PE_241_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_2_out_valid = PE_242_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_2_out_bits = PE_242_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_3_out_valid = PE_243_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_3_out_bits = PE_243_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_4_out_valid = PE_244_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_4_out_bits = PE_244_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_5_out_valid = PE_245_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_5_out_bits = PE_245_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_6_out_valid = PE_246_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_6_out_bits = PE_246_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_7_out_valid = PE_247_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_7_out_bits = PE_247_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_8_out_valid = PE_248_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_8_out_bits = PE_248_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_9_out_valid = PE_249_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_9_out_bits = PE_249_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_10_out_valid = PE_250_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_10_out_bits = PE_250_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_11_out_valid = PE_251_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_11_out_bits = PE_251_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_12_out_valid = PE_252_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_12_out_bits = PE_252_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_13_out_valid = PE_253_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_13_out_bits = PE_253_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_14_out_valid = PE_254_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_pes_14_out_bits = PE_254_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_31_io_to_mem_valid = MemController_31_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_31_io_to_mem_bits = MemController_31_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_32_io_to_pes_0_out_valid = PE_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_0_out_bits = PE_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_1_out_valid = PE_16_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_1_out_bits = PE_16_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_2_out_valid = PE_32_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_2_out_bits = PE_32_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_3_out_valid = PE_48_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_3_out_bits = PE_48_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_4_out_valid = PE_64_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_4_out_bits = PE_64_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_5_out_valid = PE_80_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_5_out_bits = PE_80_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_6_out_valid = PE_96_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_6_out_bits = PE_96_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_7_out_valid = PE_112_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_7_out_bits = PE_112_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_8_out_valid = PE_128_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_8_out_bits = PE_128_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_9_out_valid = PE_144_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_9_out_bits = PE_144_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_10_out_valid = PE_160_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_10_out_bits = PE_160_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_11_out_valid = PE_176_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_11_out_bits = PE_176_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_12_out_valid = PE_192_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_12_out_bits = PE_192_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_13_out_valid = PE_208_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_13_out_bits = PE_208_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_14_out_valid = PE_224_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_pes_14_out_bits = PE_224_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_32_io_to_mem_valid = MemController_32_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_32_io_to_mem_bits = MemController_32_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_33_io_to_pes_0_out_valid = PE_1_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_0_out_bits = PE_1_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_1_out_valid = PE_17_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_1_out_bits = PE_17_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_2_out_valid = PE_33_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_2_out_bits = PE_33_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_3_out_valid = PE_49_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_3_out_bits = PE_49_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_4_out_valid = PE_65_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_4_out_bits = PE_65_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_5_out_valid = PE_81_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_5_out_bits = PE_81_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_6_out_valid = PE_97_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_6_out_bits = PE_97_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_7_out_valid = PE_113_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_7_out_bits = PE_113_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_8_out_valid = PE_129_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_8_out_bits = PE_129_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_9_out_valid = PE_145_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_9_out_bits = PE_145_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_10_out_valid = PE_161_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_10_out_bits = PE_161_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_11_out_valid = PE_177_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_11_out_bits = PE_177_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_12_out_valid = PE_193_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_12_out_bits = PE_193_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_13_out_valid = PE_209_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_13_out_bits = PE_209_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_14_out_valid = PE_225_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_pes_14_out_bits = PE_225_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_33_io_to_mem_valid = MemController_33_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_33_io_to_mem_bits = MemController_33_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_34_io_to_pes_0_out_valid = PE_2_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_0_out_bits = PE_2_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_1_out_valid = PE_18_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_1_out_bits = PE_18_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_2_out_valid = PE_34_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_2_out_bits = PE_34_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_3_out_valid = PE_50_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_3_out_bits = PE_50_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_4_out_valid = PE_66_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_4_out_bits = PE_66_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_5_out_valid = PE_82_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_5_out_bits = PE_82_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_6_out_valid = PE_98_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_6_out_bits = PE_98_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_7_out_valid = PE_114_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_7_out_bits = PE_114_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_8_out_valid = PE_130_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_8_out_bits = PE_130_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_9_out_valid = PE_146_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_9_out_bits = PE_146_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_10_out_valid = PE_162_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_10_out_bits = PE_162_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_11_out_valid = PE_178_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_11_out_bits = PE_178_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_12_out_valid = PE_194_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_12_out_bits = PE_194_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_13_out_valid = PE_210_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_13_out_bits = PE_210_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_14_out_valid = PE_226_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_pes_14_out_bits = PE_226_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_34_io_to_mem_valid = MemController_34_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_34_io_to_mem_bits = MemController_34_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_35_io_to_pes_0_out_valid = PE_3_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_0_out_bits = PE_3_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_1_out_valid = PE_19_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_1_out_bits = PE_19_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_2_out_valid = PE_35_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_2_out_bits = PE_35_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_3_out_valid = PE_51_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_3_out_bits = PE_51_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_4_out_valid = PE_67_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_4_out_bits = PE_67_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_5_out_valid = PE_83_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_5_out_bits = PE_83_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_6_out_valid = PE_99_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_6_out_bits = PE_99_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_7_out_valid = PE_115_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_7_out_bits = PE_115_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_8_out_valid = PE_131_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_8_out_bits = PE_131_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_9_out_valid = PE_147_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_9_out_bits = PE_147_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_10_out_valid = PE_163_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_10_out_bits = PE_163_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_11_out_valid = PE_179_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_11_out_bits = PE_179_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_12_out_valid = PE_195_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_12_out_bits = PE_195_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_13_out_valid = PE_211_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_13_out_bits = PE_211_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_14_out_valid = PE_227_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_pes_14_out_bits = PE_227_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_35_io_to_mem_valid = MemController_35_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_35_io_to_mem_bits = MemController_35_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_36_io_to_pes_0_out_valid = PE_4_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_0_out_bits = PE_4_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_1_out_valid = PE_20_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_1_out_bits = PE_20_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_2_out_valid = PE_36_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_2_out_bits = PE_36_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_3_out_valid = PE_52_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_3_out_bits = PE_52_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_4_out_valid = PE_68_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_4_out_bits = PE_68_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_5_out_valid = PE_84_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_5_out_bits = PE_84_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_6_out_valid = PE_100_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_6_out_bits = PE_100_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_7_out_valid = PE_116_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_7_out_bits = PE_116_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_8_out_valid = PE_132_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_8_out_bits = PE_132_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_9_out_valid = PE_148_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_9_out_bits = PE_148_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_10_out_valid = PE_164_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_10_out_bits = PE_164_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_11_out_valid = PE_180_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_11_out_bits = PE_180_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_12_out_valid = PE_196_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_12_out_bits = PE_196_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_13_out_valid = PE_212_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_13_out_bits = PE_212_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_14_out_valid = PE_228_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_pes_14_out_bits = PE_228_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_36_io_to_mem_valid = MemController_36_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_36_io_to_mem_bits = MemController_36_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_37_io_to_pes_0_out_valid = PE_5_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_0_out_bits = PE_5_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_1_out_valid = PE_21_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_1_out_bits = PE_21_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_2_out_valid = PE_37_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_2_out_bits = PE_37_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_3_out_valid = PE_53_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_3_out_bits = PE_53_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_4_out_valid = PE_69_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_4_out_bits = PE_69_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_5_out_valid = PE_85_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_5_out_bits = PE_85_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_6_out_valid = PE_101_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_6_out_bits = PE_101_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_7_out_valid = PE_117_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_7_out_bits = PE_117_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_8_out_valid = PE_133_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_8_out_bits = PE_133_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_9_out_valid = PE_149_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_9_out_bits = PE_149_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_10_out_valid = PE_165_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_10_out_bits = PE_165_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_11_out_valid = PE_181_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_11_out_bits = PE_181_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_12_out_valid = PE_197_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_12_out_bits = PE_197_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_13_out_valid = PE_213_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_13_out_bits = PE_213_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_14_out_valid = PE_229_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_pes_14_out_bits = PE_229_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_37_io_to_mem_valid = MemController_37_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_37_io_to_mem_bits = MemController_37_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_38_io_to_pes_0_out_valid = PE_6_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_0_out_bits = PE_6_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_1_out_valid = PE_22_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_1_out_bits = PE_22_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_2_out_valid = PE_38_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_2_out_bits = PE_38_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_3_out_valid = PE_54_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_3_out_bits = PE_54_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_4_out_valid = PE_70_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_4_out_bits = PE_70_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_5_out_valid = PE_86_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_5_out_bits = PE_86_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_6_out_valid = PE_102_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_6_out_bits = PE_102_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_7_out_valid = PE_118_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_7_out_bits = PE_118_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_8_out_valid = PE_134_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_8_out_bits = PE_134_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_9_out_valid = PE_150_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_9_out_bits = PE_150_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_10_out_valid = PE_166_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_10_out_bits = PE_166_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_11_out_valid = PE_182_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_11_out_bits = PE_182_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_12_out_valid = PE_198_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_12_out_bits = PE_198_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_13_out_valid = PE_214_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_13_out_bits = PE_214_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_14_out_valid = PE_230_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_pes_14_out_bits = PE_230_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_38_io_to_mem_valid = MemController_38_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_38_io_to_mem_bits = MemController_38_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_39_io_to_pes_0_out_valid = PE_7_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_0_out_bits = PE_7_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_1_out_valid = PE_23_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_1_out_bits = PE_23_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_2_out_valid = PE_39_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_2_out_bits = PE_39_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_3_out_valid = PE_55_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_3_out_bits = PE_55_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_4_out_valid = PE_71_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_4_out_bits = PE_71_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_5_out_valid = PE_87_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_5_out_bits = PE_87_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_6_out_valid = PE_103_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_6_out_bits = PE_103_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_7_out_valid = PE_119_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_7_out_bits = PE_119_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_8_out_valid = PE_135_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_8_out_bits = PE_135_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_9_out_valid = PE_151_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_9_out_bits = PE_151_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_10_out_valid = PE_167_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_10_out_bits = PE_167_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_11_out_valid = PE_183_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_11_out_bits = PE_183_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_12_out_valid = PE_199_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_12_out_bits = PE_199_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_13_out_valid = PE_215_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_13_out_bits = PE_215_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_14_out_valid = PE_231_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_pes_14_out_bits = PE_231_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_39_io_to_mem_valid = MemController_39_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_39_io_to_mem_bits = MemController_39_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_40_io_to_pes_0_out_valid = PE_8_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_0_out_bits = PE_8_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_1_out_valid = PE_24_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_1_out_bits = PE_24_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_2_out_valid = PE_40_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_2_out_bits = PE_40_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_3_out_valid = PE_56_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_3_out_bits = PE_56_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_4_out_valid = PE_72_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_4_out_bits = PE_72_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_5_out_valid = PE_88_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_5_out_bits = PE_88_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_6_out_valid = PE_104_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_6_out_bits = PE_104_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_7_out_valid = PE_120_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_7_out_bits = PE_120_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_8_out_valid = PE_136_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_8_out_bits = PE_136_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_9_out_valid = PE_152_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_9_out_bits = PE_152_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_10_out_valid = PE_168_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_10_out_bits = PE_168_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_11_out_valid = PE_184_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_11_out_bits = PE_184_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_12_out_valid = PE_200_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_12_out_bits = PE_200_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_13_out_valid = PE_216_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_13_out_bits = PE_216_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_14_out_valid = PE_232_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_pes_14_out_bits = PE_232_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_40_io_to_mem_valid = MemController_40_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_40_io_to_mem_bits = MemController_40_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_41_io_to_pes_0_out_valid = PE_9_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_0_out_bits = PE_9_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_1_out_valid = PE_25_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_1_out_bits = PE_25_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_2_out_valid = PE_41_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_2_out_bits = PE_41_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_3_out_valid = PE_57_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_3_out_bits = PE_57_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_4_out_valid = PE_73_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_4_out_bits = PE_73_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_5_out_valid = PE_89_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_5_out_bits = PE_89_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_6_out_valid = PE_105_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_6_out_bits = PE_105_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_7_out_valid = PE_121_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_7_out_bits = PE_121_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_8_out_valid = PE_137_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_8_out_bits = PE_137_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_9_out_valid = PE_153_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_9_out_bits = PE_153_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_10_out_valid = PE_169_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_10_out_bits = PE_169_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_11_out_valid = PE_185_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_11_out_bits = PE_185_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_12_out_valid = PE_201_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_12_out_bits = PE_201_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_13_out_valid = PE_217_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_13_out_bits = PE_217_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_14_out_valid = PE_233_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_pes_14_out_bits = PE_233_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_41_io_to_mem_valid = MemController_41_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_41_io_to_mem_bits = MemController_41_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_42_io_to_pes_0_out_valid = PE_10_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_0_out_bits = PE_10_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_1_out_valid = PE_26_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_1_out_bits = PE_26_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_2_out_valid = PE_42_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_2_out_bits = PE_42_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_3_out_valid = PE_58_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_3_out_bits = PE_58_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_4_out_valid = PE_74_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_4_out_bits = PE_74_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_5_out_valid = PE_90_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_5_out_bits = PE_90_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_6_out_valid = PE_106_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_6_out_bits = PE_106_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_7_out_valid = PE_122_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_7_out_bits = PE_122_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_8_out_valid = PE_138_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_8_out_bits = PE_138_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_9_out_valid = PE_154_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_9_out_bits = PE_154_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_10_out_valid = PE_170_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_10_out_bits = PE_170_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_11_out_valid = PE_186_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_11_out_bits = PE_186_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_12_out_valid = PE_202_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_12_out_bits = PE_202_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_13_out_valid = PE_218_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_13_out_bits = PE_218_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_14_out_valid = PE_234_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_pes_14_out_bits = PE_234_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_42_io_to_mem_valid = MemController_42_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_42_io_to_mem_bits = MemController_42_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_43_io_to_pes_0_out_valid = PE_11_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_0_out_bits = PE_11_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_1_out_valid = PE_27_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_1_out_bits = PE_27_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_2_out_valid = PE_43_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_2_out_bits = PE_43_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_3_out_valid = PE_59_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_3_out_bits = PE_59_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_4_out_valid = PE_75_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_4_out_bits = PE_75_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_5_out_valid = PE_91_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_5_out_bits = PE_91_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_6_out_valid = PE_107_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_6_out_bits = PE_107_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_7_out_valid = PE_123_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_7_out_bits = PE_123_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_8_out_valid = PE_139_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_8_out_bits = PE_139_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_9_out_valid = PE_155_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_9_out_bits = PE_155_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_10_out_valid = PE_171_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_10_out_bits = PE_171_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_11_out_valid = PE_187_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_11_out_bits = PE_187_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_12_out_valid = PE_203_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_12_out_bits = PE_203_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_13_out_valid = PE_219_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_13_out_bits = PE_219_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_14_out_valid = PE_235_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_pes_14_out_bits = PE_235_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_43_io_to_mem_valid = MemController_43_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_43_io_to_mem_bits = MemController_43_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_44_io_to_pes_0_out_valid = PE_12_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_0_out_bits = PE_12_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_1_out_valid = PE_28_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_1_out_bits = PE_28_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_2_out_valid = PE_44_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_2_out_bits = PE_44_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_3_out_valid = PE_60_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_3_out_bits = PE_60_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_4_out_valid = PE_76_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_4_out_bits = PE_76_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_5_out_valid = PE_92_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_5_out_bits = PE_92_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_6_out_valid = PE_108_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_6_out_bits = PE_108_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_7_out_valid = PE_124_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_7_out_bits = PE_124_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_8_out_valid = PE_140_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_8_out_bits = PE_140_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_9_out_valid = PE_156_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_9_out_bits = PE_156_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_10_out_valid = PE_172_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_10_out_bits = PE_172_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_11_out_valid = PE_188_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_11_out_bits = PE_188_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_12_out_valid = PE_204_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_12_out_bits = PE_204_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_13_out_valid = PE_220_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_13_out_bits = PE_220_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_14_out_valid = PE_236_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_pes_14_out_bits = PE_236_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_44_io_to_mem_valid = MemController_44_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_44_io_to_mem_bits = MemController_44_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_45_io_to_pes_0_out_valid = PE_13_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_0_out_bits = PE_13_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_1_out_valid = PE_29_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_1_out_bits = PE_29_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_2_out_valid = PE_45_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_2_out_bits = PE_45_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_3_out_valid = PE_61_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_3_out_bits = PE_61_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_4_out_valid = PE_77_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_4_out_bits = PE_77_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_5_out_valid = PE_93_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_5_out_bits = PE_93_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_6_out_valid = PE_109_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_6_out_bits = PE_109_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_7_out_valid = PE_125_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_7_out_bits = PE_125_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_8_out_valid = PE_141_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_8_out_bits = PE_141_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_9_out_valid = PE_157_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_9_out_bits = PE_157_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_10_out_valid = PE_173_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_10_out_bits = PE_173_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_11_out_valid = PE_189_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_11_out_bits = PE_189_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_12_out_valid = PE_205_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_12_out_bits = PE_205_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_13_out_valid = PE_221_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_13_out_bits = PE_221_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_14_out_valid = PE_237_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_pes_14_out_bits = PE_237_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_45_io_to_mem_valid = MemController_45_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_45_io_to_mem_bits = MemController_45_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_46_io_to_pes_0_out_valid = PE_14_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_0_out_bits = PE_14_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_1_out_valid = PE_30_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_1_out_bits = PE_30_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_2_out_valid = PE_46_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_2_out_bits = PE_46_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_3_out_valid = PE_62_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_3_out_bits = PE_62_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_4_out_valid = PE_78_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_4_out_bits = PE_78_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_5_out_valid = PE_94_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_5_out_bits = PE_94_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_6_out_valid = PE_110_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_6_out_bits = PE_110_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_7_out_valid = PE_126_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_7_out_bits = PE_126_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_8_out_valid = PE_142_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_8_out_bits = PE_142_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_9_out_valid = PE_158_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_9_out_bits = PE_158_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_10_out_valid = PE_174_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_10_out_bits = PE_174_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_11_out_valid = PE_190_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_11_out_bits = PE_190_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_12_out_valid = PE_206_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_12_out_bits = PE_206_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_13_out_valid = PE_222_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_13_out_bits = PE_222_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_14_out_valid = PE_238_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_pes_14_out_bits = PE_238_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_46_io_to_mem_valid = MemController_46_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_46_io_to_mem_bits = MemController_46_io_rd_data_bits; // @[pearray.scala 255:29]
  assign PENetwork_47_io_to_pes_0_out_valid = PE_15_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_0_out_bits = PE_15_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_1_out_valid = PE_31_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_1_out_bits = PE_31_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_2_out_valid = PE_47_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_2_out_bits = PE_47_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_3_out_valid = PE_63_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_3_out_bits = PE_63_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_4_out_valid = PE_79_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_4_out_bits = PE_79_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_5_out_valid = PE_95_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_5_out_bits = PE_95_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_6_out_valid = PE_111_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_6_out_bits = PE_111_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_7_out_valid = PE_127_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_7_out_bits = PE_127_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_8_out_valid = PE_143_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_8_out_bits = PE_143_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_9_out_valid = PE_159_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_9_out_bits = PE_159_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_10_out_valid = PE_175_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_10_out_bits = PE_175_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_11_out_valid = PE_191_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_11_out_bits = PE_191_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_12_out_valid = PE_207_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_12_out_bits = PE_207_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_13_out_valid = PE_223_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_13_out_bits = PE_223_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_14_out_valid = PE_239_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_pes_14_out_bits = PE_239_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_47_io_to_mem_valid = MemController_47_io_rd_data_valid; // @[pearray.scala 255:29]
  assign PENetwork_47_io_to_mem_bits = MemController_47_io_rd_data_bits; // @[pearray.scala 255:29]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_io_wr_valid = PENetwork_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_io_wr_data_valid = PENetwork_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_io_wr_data_bits = PENetwork_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_1_clock = clock;
  assign MemController_1_reset = reset;
  assign MemController_1_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_1_io_wr_valid = PENetwork_1_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_1_io_wr_data_valid = PENetwork_1_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_1_io_wr_data_bits = PENetwork_1_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_2_clock = clock;
  assign MemController_2_reset = reset;
  assign MemController_2_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_2_io_wr_valid = PENetwork_2_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_2_io_wr_data_valid = PENetwork_2_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_2_io_wr_data_bits = PENetwork_2_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_3_clock = clock;
  assign MemController_3_reset = reset;
  assign MemController_3_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_3_io_wr_valid = PENetwork_3_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_3_io_wr_data_valid = PENetwork_3_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_3_io_wr_data_bits = PENetwork_3_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_4_clock = clock;
  assign MemController_4_reset = reset;
  assign MemController_4_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_4_io_wr_valid = PENetwork_4_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_4_io_wr_data_valid = PENetwork_4_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_4_io_wr_data_bits = PENetwork_4_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_5_clock = clock;
  assign MemController_5_reset = reset;
  assign MemController_5_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_5_io_wr_valid = PENetwork_5_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_5_io_wr_data_valid = PENetwork_5_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_5_io_wr_data_bits = PENetwork_5_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_6_clock = clock;
  assign MemController_6_reset = reset;
  assign MemController_6_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_6_io_wr_valid = PENetwork_6_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_6_io_wr_data_valid = PENetwork_6_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_6_io_wr_data_bits = PENetwork_6_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_7_clock = clock;
  assign MemController_7_reset = reset;
  assign MemController_7_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_7_io_wr_valid = PENetwork_7_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_7_io_wr_data_valid = PENetwork_7_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_7_io_wr_data_bits = PENetwork_7_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_8_clock = clock;
  assign MemController_8_reset = reset;
  assign MemController_8_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_8_io_wr_valid = PENetwork_8_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_8_io_wr_data_valid = PENetwork_8_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_8_io_wr_data_bits = PENetwork_8_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_9_clock = clock;
  assign MemController_9_reset = reset;
  assign MemController_9_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_9_io_wr_valid = PENetwork_9_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_9_io_wr_data_valid = PENetwork_9_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_9_io_wr_data_bits = PENetwork_9_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_10_clock = clock;
  assign MemController_10_reset = reset;
  assign MemController_10_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_10_io_wr_valid = PENetwork_10_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_10_io_wr_data_valid = PENetwork_10_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_10_io_wr_data_bits = PENetwork_10_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_11_clock = clock;
  assign MemController_11_reset = reset;
  assign MemController_11_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_11_io_wr_valid = PENetwork_11_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_11_io_wr_data_valid = PENetwork_11_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_11_io_wr_data_bits = PENetwork_11_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_12_clock = clock;
  assign MemController_12_reset = reset;
  assign MemController_12_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_12_io_wr_valid = PENetwork_12_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_12_io_wr_data_valid = PENetwork_12_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_12_io_wr_data_bits = PENetwork_12_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_13_clock = clock;
  assign MemController_13_reset = reset;
  assign MemController_13_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_13_io_wr_valid = PENetwork_13_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_13_io_wr_data_valid = PENetwork_13_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_13_io_wr_data_bits = PENetwork_13_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_14_clock = clock;
  assign MemController_14_reset = reset;
  assign MemController_14_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_14_io_wr_valid = PENetwork_14_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_14_io_wr_data_valid = PENetwork_14_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_14_io_wr_data_bits = PENetwork_14_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_15_clock = clock;
  assign MemController_15_reset = reset;
  assign MemController_15_io_rd_valid = io_out_valid; // @[pearray.scala 259:28]
  assign MemController_15_io_wr_valid = PENetwork_15_io_to_mem_valid; // @[pearray.scala 258:28]
  assign MemController_15_io_wr_data_valid = PENetwork_15_io_to_mem_valid; // @[pearray.scala 260:27]
  assign MemController_15_io_wr_data_bits = PENetwork_15_io_to_mem_bits; // @[pearray.scala 260:27]
  assign MemController_16_clock = clock;
  assign MemController_16_reset = reset;
  assign MemController_16_io_rd_valid = _T_2575_2; // @[pearray.scala 252:30]
  assign MemController_16_io_wr_valid = io_data_1_in_0_valid; // @[pearray.scala 253:28]
  assign MemController_16_io_wr_data_valid = io_data_1_in_0_bits_valid; // @[pearray.scala 254:27]
  assign MemController_16_io_wr_data_bits = io_data_1_in_0_bits_bits; // @[pearray.scala 254:27]
  assign MemController_17_clock = clock;
  assign MemController_17_reset = reset;
  assign MemController_17_io_rd_valid = _T_2584_2; // @[pearray.scala 252:30]
  assign MemController_17_io_wr_valid = io_data_1_in_1_valid; // @[pearray.scala 253:28]
  assign MemController_17_io_wr_data_valid = io_data_1_in_1_bits_valid; // @[pearray.scala 254:27]
  assign MemController_17_io_wr_data_bits = io_data_1_in_1_bits_bits; // @[pearray.scala 254:27]
  assign MemController_18_clock = clock;
  assign MemController_18_reset = reset;
  assign MemController_18_io_rd_valid = _T_2593_2; // @[pearray.scala 252:30]
  assign MemController_18_io_wr_valid = io_data_1_in_2_valid; // @[pearray.scala 253:28]
  assign MemController_18_io_wr_data_valid = io_data_1_in_2_bits_valid; // @[pearray.scala 254:27]
  assign MemController_18_io_wr_data_bits = io_data_1_in_2_bits_bits; // @[pearray.scala 254:27]
  assign MemController_19_clock = clock;
  assign MemController_19_reset = reset;
  assign MemController_19_io_rd_valid = _T_2602_2; // @[pearray.scala 252:30]
  assign MemController_19_io_wr_valid = io_data_1_in_3_valid; // @[pearray.scala 253:28]
  assign MemController_19_io_wr_data_valid = io_data_1_in_3_bits_valid; // @[pearray.scala 254:27]
  assign MemController_19_io_wr_data_bits = io_data_1_in_3_bits_bits; // @[pearray.scala 254:27]
  assign MemController_20_clock = clock;
  assign MemController_20_reset = reset;
  assign MemController_20_io_rd_valid = _T_2611_2; // @[pearray.scala 252:30]
  assign MemController_20_io_wr_valid = io_data_1_in_4_valid; // @[pearray.scala 253:28]
  assign MemController_20_io_wr_data_valid = io_data_1_in_4_bits_valid; // @[pearray.scala 254:27]
  assign MemController_20_io_wr_data_bits = io_data_1_in_4_bits_bits; // @[pearray.scala 254:27]
  assign MemController_21_clock = clock;
  assign MemController_21_reset = reset;
  assign MemController_21_io_rd_valid = _T_2620_2; // @[pearray.scala 252:30]
  assign MemController_21_io_wr_valid = io_data_1_in_5_valid; // @[pearray.scala 253:28]
  assign MemController_21_io_wr_data_valid = io_data_1_in_5_bits_valid; // @[pearray.scala 254:27]
  assign MemController_21_io_wr_data_bits = io_data_1_in_5_bits_bits; // @[pearray.scala 254:27]
  assign MemController_22_clock = clock;
  assign MemController_22_reset = reset;
  assign MemController_22_io_rd_valid = _T_2629_2; // @[pearray.scala 252:30]
  assign MemController_22_io_wr_valid = io_data_1_in_6_valid; // @[pearray.scala 253:28]
  assign MemController_22_io_wr_data_valid = io_data_1_in_6_bits_valid; // @[pearray.scala 254:27]
  assign MemController_22_io_wr_data_bits = io_data_1_in_6_bits_bits; // @[pearray.scala 254:27]
  assign MemController_23_clock = clock;
  assign MemController_23_reset = reset;
  assign MemController_23_io_rd_valid = _T_2638_2; // @[pearray.scala 252:30]
  assign MemController_23_io_wr_valid = io_data_1_in_7_valid; // @[pearray.scala 253:28]
  assign MemController_23_io_wr_data_valid = io_data_1_in_7_bits_valid; // @[pearray.scala 254:27]
  assign MemController_23_io_wr_data_bits = io_data_1_in_7_bits_bits; // @[pearray.scala 254:27]
  assign MemController_24_clock = clock;
  assign MemController_24_reset = reset;
  assign MemController_24_io_rd_valid = _T_2647_2; // @[pearray.scala 252:30]
  assign MemController_24_io_wr_valid = io_data_1_in_8_valid; // @[pearray.scala 253:28]
  assign MemController_24_io_wr_data_valid = io_data_1_in_8_bits_valid; // @[pearray.scala 254:27]
  assign MemController_24_io_wr_data_bits = io_data_1_in_8_bits_bits; // @[pearray.scala 254:27]
  assign MemController_25_clock = clock;
  assign MemController_25_reset = reset;
  assign MemController_25_io_rd_valid = _T_2656_2; // @[pearray.scala 252:30]
  assign MemController_25_io_wr_valid = io_data_1_in_9_valid; // @[pearray.scala 253:28]
  assign MemController_25_io_wr_data_valid = io_data_1_in_9_bits_valid; // @[pearray.scala 254:27]
  assign MemController_25_io_wr_data_bits = io_data_1_in_9_bits_bits; // @[pearray.scala 254:27]
  assign MemController_26_clock = clock;
  assign MemController_26_reset = reset;
  assign MemController_26_io_rd_valid = _T_2665_2; // @[pearray.scala 252:30]
  assign MemController_26_io_wr_valid = io_data_1_in_10_valid; // @[pearray.scala 253:28]
  assign MemController_26_io_wr_data_valid = io_data_1_in_10_bits_valid; // @[pearray.scala 254:27]
  assign MemController_26_io_wr_data_bits = io_data_1_in_10_bits_bits; // @[pearray.scala 254:27]
  assign MemController_27_clock = clock;
  assign MemController_27_reset = reset;
  assign MemController_27_io_rd_valid = _T_2674_2; // @[pearray.scala 252:30]
  assign MemController_27_io_wr_valid = io_data_1_in_11_valid; // @[pearray.scala 253:28]
  assign MemController_27_io_wr_data_valid = io_data_1_in_11_bits_valid; // @[pearray.scala 254:27]
  assign MemController_27_io_wr_data_bits = io_data_1_in_11_bits_bits; // @[pearray.scala 254:27]
  assign MemController_28_clock = clock;
  assign MemController_28_reset = reset;
  assign MemController_28_io_rd_valid = _T_2683_2; // @[pearray.scala 252:30]
  assign MemController_28_io_wr_valid = io_data_1_in_12_valid; // @[pearray.scala 253:28]
  assign MemController_28_io_wr_data_valid = io_data_1_in_12_bits_valid; // @[pearray.scala 254:27]
  assign MemController_28_io_wr_data_bits = io_data_1_in_12_bits_bits; // @[pearray.scala 254:27]
  assign MemController_29_clock = clock;
  assign MemController_29_reset = reset;
  assign MemController_29_io_rd_valid = _T_2692_2; // @[pearray.scala 252:30]
  assign MemController_29_io_wr_valid = io_data_1_in_13_valid; // @[pearray.scala 253:28]
  assign MemController_29_io_wr_data_valid = io_data_1_in_13_bits_valid; // @[pearray.scala 254:27]
  assign MemController_29_io_wr_data_bits = io_data_1_in_13_bits_bits; // @[pearray.scala 254:27]
  assign MemController_30_clock = clock;
  assign MemController_30_reset = reset;
  assign MemController_30_io_rd_valid = _T_2701_2; // @[pearray.scala 252:30]
  assign MemController_30_io_wr_valid = io_data_1_in_14_valid; // @[pearray.scala 253:28]
  assign MemController_30_io_wr_data_valid = io_data_1_in_14_bits_valid; // @[pearray.scala 254:27]
  assign MemController_30_io_wr_data_bits = io_data_1_in_14_bits_bits; // @[pearray.scala 254:27]
  assign MemController_31_clock = clock;
  assign MemController_31_reset = reset;
  assign MemController_31_io_rd_valid = _T_2710_2; // @[pearray.scala 252:30]
  assign MemController_31_io_wr_valid = io_data_1_in_15_valid; // @[pearray.scala 253:28]
  assign MemController_31_io_wr_data_valid = io_data_1_in_15_bits_valid; // @[pearray.scala 254:27]
  assign MemController_31_io_wr_data_bits = io_data_1_in_15_bits_bits; // @[pearray.scala 254:27]
  assign MemController_32_clock = clock;
  assign MemController_32_reset = reset;
  assign MemController_32_io_rd_valid = io_exec_valid; // @[pearray.scala 245:32]
  assign MemController_32_io_wr_valid = io_data_2_in_0_valid; // @[pearray.scala 253:28]
  assign MemController_32_io_wr_data_valid = io_data_2_in_0_bits_valid; // @[pearray.scala 254:27]
  assign MemController_32_io_wr_data_bits = io_data_2_in_0_bits_bits; // @[pearray.scala 254:27]
  assign MemController_33_clock = clock;
  assign MemController_33_reset = reset;
  assign MemController_33_io_rd_valid = _T_2712_11; // @[pearray.scala 243:32]
  assign MemController_33_io_wr_valid = io_data_2_in_1_valid; // @[pearray.scala 253:28]
  assign MemController_33_io_wr_data_valid = io_data_2_in_1_bits_valid; // @[pearray.scala 254:27]
  assign MemController_33_io_wr_data_bits = io_data_2_in_1_bits_bits; // @[pearray.scala 254:27]
  assign MemController_34_clock = clock;
  assign MemController_34_reset = reset;
  assign MemController_34_io_rd_valid = _T_2712_23; // @[pearray.scala 243:32]
  assign MemController_34_io_wr_valid = io_data_2_in_2_valid; // @[pearray.scala 253:28]
  assign MemController_34_io_wr_data_valid = io_data_2_in_2_bits_valid; // @[pearray.scala 254:27]
  assign MemController_34_io_wr_data_bits = io_data_2_in_2_bits_bits; // @[pearray.scala 254:27]
  assign MemController_35_clock = clock;
  assign MemController_35_reset = reset;
  assign MemController_35_io_rd_valid = _T_2712_35; // @[pearray.scala 243:32]
  assign MemController_35_io_wr_valid = io_data_2_in_3_valid; // @[pearray.scala 253:28]
  assign MemController_35_io_wr_data_valid = io_data_2_in_3_bits_valid; // @[pearray.scala 254:27]
  assign MemController_35_io_wr_data_bits = io_data_2_in_3_bits_bits; // @[pearray.scala 254:27]
  assign MemController_36_clock = clock;
  assign MemController_36_reset = reset;
  assign MemController_36_io_rd_valid = _T_2712_47; // @[pearray.scala 243:32]
  assign MemController_36_io_wr_valid = io_data_2_in_4_valid; // @[pearray.scala 253:28]
  assign MemController_36_io_wr_data_valid = io_data_2_in_4_bits_valid; // @[pearray.scala 254:27]
  assign MemController_36_io_wr_data_bits = io_data_2_in_4_bits_bits; // @[pearray.scala 254:27]
  assign MemController_37_clock = clock;
  assign MemController_37_reset = reset;
  assign MemController_37_io_rd_valid = _T_2712_59; // @[pearray.scala 243:32]
  assign MemController_37_io_wr_valid = io_data_2_in_5_valid; // @[pearray.scala 253:28]
  assign MemController_37_io_wr_data_valid = io_data_2_in_5_bits_valid; // @[pearray.scala 254:27]
  assign MemController_37_io_wr_data_bits = io_data_2_in_5_bits_bits; // @[pearray.scala 254:27]
  assign MemController_38_clock = clock;
  assign MemController_38_reset = reset;
  assign MemController_38_io_rd_valid = _T_2712_71; // @[pearray.scala 243:32]
  assign MemController_38_io_wr_valid = io_data_2_in_6_valid; // @[pearray.scala 253:28]
  assign MemController_38_io_wr_data_valid = io_data_2_in_6_bits_valid; // @[pearray.scala 254:27]
  assign MemController_38_io_wr_data_bits = io_data_2_in_6_bits_bits; // @[pearray.scala 254:27]
  assign MemController_39_clock = clock;
  assign MemController_39_reset = reset;
  assign MemController_39_io_rd_valid = _T_2712_83; // @[pearray.scala 243:32]
  assign MemController_39_io_wr_valid = io_data_2_in_7_valid; // @[pearray.scala 253:28]
  assign MemController_39_io_wr_data_valid = io_data_2_in_7_bits_valid; // @[pearray.scala 254:27]
  assign MemController_39_io_wr_data_bits = io_data_2_in_7_bits_bits; // @[pearray.scala 254:27]
  assign MemController_40_clock = clock;
  assign MemController_40_reset = reset;
  assign MemController_40_io_rd_valid = _T_2712_95; // @[pearray.scala 243:32]
  assign MemController_40_io_wr_valid = io_data_2_in_8_valid; // @[pearray.scala 253:28]
  assign MemController_40_io_wr_data_valid = io_data_2_in_8_bits_valid; // @[pearray.scala 254:27]
  assign MemController_40_io_wr_data_bits = io_data_2_in_8_bits_bits; // @[pearray.scala 254:27]
  assign MemController_41_clock = clock;
  assign MemController_41_reset = reset;
  assign MemController_41_io_rd_valid = _T_2712_107; // @[pearray.scala 243:32]
  assign MemController_41_io_wr_valid = io_data_2_in_9_valid; // @[pearray.scala 253:28]
  assign MemController_41_io_wr_data_valid = io_data_2_in_9_bits_valid; // @[pearray.scala 254:27]
  assign MemController_41_io_wr_data_bits = io_data_2_in_9_bits_bits; // @[pearray.scala 254:27]
  assign MemController_42_clock = clock;
  assign MemController_42_reset = reset;
  assign MemController_42_io_rd_valid = _T_2712_119; // @[pearray.scala 243:32]
  assign MemController_42_io_wr_valid = io_data_2_in_10_valid; // @[pearray.scala 253:28]
  assign MemController_42_io_wr_data_valid = io_data_2_in_10_bits_valid; // @[pearray.scala 254:27]
  assign MemController_42_io_wr_data_bits = io_data_2_in_10_bits_bits; // @[pearray.scala 254:27]
  assign MemController_43_clock = clock;
  assign MemController_43_reset = reset;
  assign MemController_43_io_rd_valid = _T_2712_131; // @[pearray.scala 243:32]
  assign MemController_43_io_wr_valid = io_data_2_in_11_valid; // @[pearray.scala 253:28]
  assign MemController_43_io_wr_data_valid = io_data_2_in_11_bits_valid; // @[pearray.scala 254:27]
  assign MemController_43_io_wr_data_bits = io_data_2_in_11_bits_bits; // @[pearray.scala 254:27]
  assign MemController_44_clock = clock;
  assign MemController_44_reset = reset;
  assign MemController_44_io_rd_valid = _T_2712_143; // @[pearray.scala 243:32]
  assign MemController_44_io_wr_valid = io_data_2_in_12_valid; // @[pearray.scala 253:28]
  assign MemController_44_io_wr_data_valid = io_data_2_in_12_bits_valid; // @[pearray.scala 254:27]
  assign MemController_44_io_wr_data_bits = io_data_2_in_12_bits_bits; // @[pearray.scala 254:27]
  assign MemController_45_clock = clock;
  assign MemController_45_reset = reset;
  assign MemController_45_io_rd_valid = _T_2712_155; // @[pearray.scala 243:32]
  assign MemController_45_io_wr_valid = io_data_2_in_13_valid; // @[pearray.scala 253:28]
  assign MemController_45_io_wr_data_valid = io_data_2_in_13_bits_valid; // @[pearray.scala 254:27]
  assign MemController_45_io_wr_data_bits = io_data_2_in_13_bits_bits; // @[pearray.scala 254:27]
  assign MemController_46_clock = clock;
  assign MemController_46_reset = reset;
  assign MemController_46_io_rd_valid = _T_2712_167; // @[pearray.scala 243:32]
  assign MemController_46_io_wr_valid = io_data_2_in_14_valid; // @[pearray.scala 253:28]
  assign MemController_46_io_wr_data_valid = io_data_2_in_14_bits_valid; // @[pearray.scala 254:27]
  assign MemController_46_io_wr_data_bits = io_data_2_in_14_bits_bits; // @[pearray.scala 254:27]
  assign MemController_47_clock = clock;
  assign MemController_47_reset = reset;
  assign MemController_47_io_rd_valid = _T_2712_179; // @[pearray.scala 243:32]
  assign MemController_47_io_wr_valid = io_data_2_in_15_valid; // @[pearray.scala 253:28]
  assign MemController_47_io_wr_data_valid = io_data_2_in_15_bits_valid; // @[pearray.scala 254:27]
  assign MemController_47_io_wr_data_bits = io_data_2_in_15_bits_bits; // @[pearray.scala 254:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_12_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_12_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_12_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_22_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_22_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_22_2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_22_3 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_32_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_32_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_32_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_32_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_42_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_42_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_42_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_42_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_52_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_52_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_52_2 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_52_3 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_62_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_62_1 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_62_2 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_62_3 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_72_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_72_1 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_72_2 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_72_3 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_82_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_82_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_82_2 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_82_3 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_92_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_92_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_92_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_92_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_102_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_102_1 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_102_2 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_102_3 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_112_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_112_1 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_112_2 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_112_3 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_122_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_122_1 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_122_2 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_122_3 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_132_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_132_1 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_132_2 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_132_3 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_142_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_142_1 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_142_2 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_142_3 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_152_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_152_1 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_152_2 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_152_3 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_162_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_162_1 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_162_2 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_162_3 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_172_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_172_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_172_2 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_172_3 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_182_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_182_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_182_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_182_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_192_0 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_192_1 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_192_2 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_192_3 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_202_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_202_1 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_202_2 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_202_3 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_212_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_212_1 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_212_2 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_212_3 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_222_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_222_1 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_222_2 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_222_3 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_232_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_232_1 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_232_2 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_232_3 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_242_0 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_242_1 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_242_2 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_242_3 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_252_0 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_252_1 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_252_2 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_252_3 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_262_0 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_262_1 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_262_2 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_262_3 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_272_0 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_272_1 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_272_2 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_272_3 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_282_0 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_282_1 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_282_2 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_282_3 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_292_0 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_292_1 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_292_2 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_292_3 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_302_0 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_302_1 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_302_2 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_302_3 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_312_0 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_312_1 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_312_2 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_312_3 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_322_0 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_322_1 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_322_2 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_322_3 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_332_0 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_332_1 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_332_2 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_332_3 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_342_0 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_342_1 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_342_2 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_342_3 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_352_0 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_352_1 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_352_2 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_352_3 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_362_0 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_362_1 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_362_2 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_362_3 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_372_0 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_372_1 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_372_2 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_372_3 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_382_0 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_382_1 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_382_2 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_382_3 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_392_0 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_392_1 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_392_2 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_392_3 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_402_0 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_402_1 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_402_2 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_402_3 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_412_0 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_412_1 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_412_2 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_412_3 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_422_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_422_1 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_422_2 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_422_3 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_432_0 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_432_1 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_432_2 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_432_3 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_442_0 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_442_1 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_442_2 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_442_3 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_452_0 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_452_1 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_452_2 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_452_3 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_462_0 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_462_1 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_462_2 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_462_3 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_472_0 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_472_1 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_472_2 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_472_3 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_482_0 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_482_1 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_482_2 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_482_3 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_492_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_492_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_492_2 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_492_3 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_502_0 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_502_1 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_502_2 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_502_3 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_512_0 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_512_1 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_512_2 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_512_3 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_522_0 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_522_1 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_522_2 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_522_3 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_532_0 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_532_1 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_532_2 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_532_3 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_542_0 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_542_1 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_542_2 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_542_3 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_552_0 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_552_1 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_552_2 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_552_3 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_562_0 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_562_1 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_562_2 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_562_3 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_572_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_572_1 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_572_2 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_572_3 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_582_0 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_582_1 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_582_2 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_582_3 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_592_0 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_592_1 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_592_2 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_592_3 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_602_0 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_602_1 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_602_2 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_602_3 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_612_0 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_612_1 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_612_2 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_612_3 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_622_0 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_622_1 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_622_2 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_622_3 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_632_0 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_632_1 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_632_2 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_632_3 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_642_0 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_642_1 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_642_2 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_642_3 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_652_0 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_652_1 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_652_2 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_652_3 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_662_0 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_662_1 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_662_2 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_662_3 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_672_0 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_672_1 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_672_2 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_672_3 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_682_0 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_682_1 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_682_2 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_682_3 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_692_0 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_692_1 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_692_2 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_692_3 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_702_0 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_702_1 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_702_2 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_702_3 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_712_0 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_712_1 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_712_2 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_712_3 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_722_0 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_722_1 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_722_2 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_722_3 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_732_0 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_732_1 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_732_2 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_732_3 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_742_0 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_742_1 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_742_2 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_742_3 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_752_0 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_752_1 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_752_2 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_752_3 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_762_0 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_762_1 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_762_2 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_762_3 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_772_0 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_772_1 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_772_2 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_772_3 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_782_0 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_782_1 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_782_2 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_782_3 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_792_0 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_792_1 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_792_2 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_792_3 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_802_0 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_802_1 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_802_2 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_802_3 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_812_0 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_812_1 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_812_2 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_812_3 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_822_0 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_822_1 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_822_2 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_822_3 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_832_0 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_832_1 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_832_2 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_832_3 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_842_0 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_842_1 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_842_2 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_842_3 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_852_0 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_852_1 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_852_2 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_852_3 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_862_0 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_862_1 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_862_2 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_862_3 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_872_0 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_872_1 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_872_2 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_872_3 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_882_0 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_882_1 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_882_2 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_882_3 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_892_0 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_892_1 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_892_2 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_892_3 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_902_0 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_902_1 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_902_2 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_902_3 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_912_0 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_912_1 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_912_2 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_912_3 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_922_0 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_922_1 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_922_2 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_922_3 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_932_0 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_932_1 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_932_2 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_932_3 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_942_0 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_942_1 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_942_2 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_942_3 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_952_0 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_952_1 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_952_2 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_952_3 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_962_0 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_962_1 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_962_2 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_962_3 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_972_0 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_972_1 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_972_2 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_972_3 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_982_0 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_982_1 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_982_2 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_982_3 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_992_0 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_992_1 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_992_2 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_992_3 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_1002_0 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_1002_1 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_1002_2 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_1002_3 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_1012_0 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_1012_1 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_1012_2 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_1012_3 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_1022_0 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_1022_1 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_1022_2 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_1022_3 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_1032_0 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_1032_1 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_1032_2 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_1032_3 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_1042_0 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_1042_1 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_1042_2 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_1042_3 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_1052_0 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_1052_1 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_1052_2 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_1052_3 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_1062_0 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_1062_1 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_1062_2 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_1062_3 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_1072_0 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_1072_1 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_1072_2 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_1072_3 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_1082_0 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_1082_1 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_1082_2 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_1082_3 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_1092_0 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_1092_1 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_1092_2 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_1092_3 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_1102_0 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_1102_1 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_1102_2 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_1102_3 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_1112_0 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_1112_1 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_1112_2 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_1112_3 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_1122_0 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_1122_1 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_1122_2 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_1122_3 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_1132_0 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_1132_1 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_1132_2 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_1132_3 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_1142_0 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_1142_1 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_1142_2 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_1142_3 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_1152_0 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_1152_1 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_1152_2 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_1152_3 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_1162_0 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_1162_1 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_1162_2 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_1162_3 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_1172_0 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_1172_1 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_1172_2 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_1172_3 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_1182_0 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_1182_1 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_1182_2 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_1182_3 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_1192_0 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_1192_1 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_1192_2 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_1192_3 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_1202_0 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_1202_1 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_1202_2 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_1202_3 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_1212_0 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_1212_1 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_1212_2 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_1212_3 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_1222_0 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_1222_1 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_1222_2 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_1222_3 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_1232_0 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_1232_1 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_1232_2 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_1232_3 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_1242_0 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_1242_1 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_1242_2 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_1242_3 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_1252_0 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_1252_1 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_1252_2 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_1252_3 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_1262_0 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_1262_1 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_1262_2 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_1262_3 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_1272_0 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_1272_1 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_1272_2 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_1272_3 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_1282_0 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_1282_1 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_1282_2 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_1282_3 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_1292_0 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_1292_1 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_1292_2 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_1292_3 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_1302_0 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_1302_1 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_1302_2 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_1302_3 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_1312_0 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_1312_1 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_1312_2 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_1312_3 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_1322_0 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_1322_1 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_1322_2 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_1322_3 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_1332_0 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_1332_1 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_1332_2 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_1332_3 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_1342_0 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_1342_1 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_1342_2 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_1342_3 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_1352_0 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_1352_1 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_1352_2 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_1352_3 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_1362_0 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_1362_1 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_1362_2 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_1362_3 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_1372_0 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_1372_1 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_1372_2 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_1372_3 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_1382_0 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_1382_1 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_1382_2 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_1382_3 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_1392_0 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_1392_1 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_1392_2 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_1392_3 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_1402_0 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_1402_1 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_1402_2 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_1402_3 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_1412_0 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_1412_1 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_1412_2 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_1412_3 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_1422_0 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_1422_1 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_1422_2 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_1422_3 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_1432_0 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_1432_1 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_1432_2 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_1432_3 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_1442_0 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_1442_1 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_1442_2 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_1442_3 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_1452_0 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_1452_1 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_1452_2 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_1452_3 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_1462_0 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_1462_1 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_1462_2 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_1462_3 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_1472_0 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_1472_1 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_1472_2 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_1472_3 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_1482_0 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_1482_1 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_1482_2 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_1482_3 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_1492_0 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_1492_1 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_1492_2 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_1492_3 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_1502_0 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_1502_1 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_1502_2 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_1502_3 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_1512_0 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_1512_1 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_1512_2 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_1512_3 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_1522_0 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_1522_1 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_1522_2 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_1522_3 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_1532_0 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_1532_1 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_1532_2 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_1532_3 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_1542_0 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_1542_1 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_1542_2 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_1542_3 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_1552_0 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_1552_1 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_1552_2 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_1552_3 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_1562_0 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_1562_1 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_1562_2 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_1562_3 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_1572_0 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_1572_1 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_1572_2 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_1572_3 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_1582_0 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_1582_1 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_1582_2 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_1582_3 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_1592_0 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_1592_1 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_1592_2 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_1592_3 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_1602_0 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_1602_1 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_1602_2 = _RAND_638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_1602_3 = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_1612_0 = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_1612_1 = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_1612_2 = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_1612_3 = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_1622_0 = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_1622_1 = _RAND_645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_1622_2 = _RAND_646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_1622_3 = _RAND_647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_1632_0 = _RAND_648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_1632_1 = _RAND_649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_1632_2 = _RAND_650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_1632_3 = _RAND_651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_1642_0 = _RAND_652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_1642_1 = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_1642_2 = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_1642_3 = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_1652_0 = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_1652_1 = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_1652_2 = _RAND_658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_1652_3 = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_1662_0 = _RAND_660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_1662_1 = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_1662_2 = _RAND_662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_1662_3 = _RAND_663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_1672_0 = _RAND_664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_1672_1 = _RAND_665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_1672_2 = _RAND_666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_1672_3 = _RAND_667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_1682_0 = _RAND_668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_1682_1 = _RAND_669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_1682_2 = _RAND_670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_1682_3 = _RAND_671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_1692_0 = _RAND_672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_1692_1 = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_1692_2 = _RAND_674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_1692_3 = _RAND_675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_1702_0 = _RAND_676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_1702_1 = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_1702_2 = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_1702_3 = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_1712_0 = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_1712_1 = _RAND_681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_1712_2 = _RAND_682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_1712_3 = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_1722_0 = _RAND_684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_1722_1 = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_1722_2 = _RAND_686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_1722_3 = _RAND_687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_1732_0 = _RAND_688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_1732_1 = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_1732_2 = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_1732_3 = _RAND_691[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_1742_0 = _RAND_692[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_1742_1 = _RAND_693[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_1742_2 = _RAND_694[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_1742_3 = _RAND_695[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_1752_0 = _RAND_696[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_1752_1 = _RAND_697[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_1752_2 = _RAND_698[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_1752_3 = _RAND_699[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_1762_0 = _RAND_700[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_1762_1 = _RAND_701[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_1762_2 = _RAND_702[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_1762_3 = _RAND_703[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_1772_0 = _RAND_704[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_1772_1 = _RAND_705[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_1772_2 = _RAND_706[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_1772_3 = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_1782_0 = _RAND_708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_1782_1 = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_1782_2 = _RAND_710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_1782_3 = _RAND_711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_1792_0 = _RAND_712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_1792_1 = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_1792_2 = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_1792_3 = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_1802_0 = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_1802_1 = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_1802_2 = _RAND_718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_1802_3 = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_1812_0 = _RAND_720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_1812_1 = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_1812_2 = _RAND_722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_1812_3 = _RAND_723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_1822_0 = _RAND_724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_1822_1 = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_1822_2 = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_1822_3 = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_1832_0 = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_1832_1 = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_1832_2 = _RAND_730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_1832_3 = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_1842_0 = _RAND_732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_1842_1 = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_1842_2 = _RAND_734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_1842_3 = _RAND_735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_1852_0 = _RAND_736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_1852_1 = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_1852_2 = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_1852_3 = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_1862_0 = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_1862_1 = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_1862_2 = _RAND_742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_1862_3 = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_1872_0 = _RAND_744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_1872_1 = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_1872_2 = _RAND_746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_1872_3 = _RAND_747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_1882_0 = _RAND_748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_1882_1 = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_1882_2 = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_1882_3 = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_1892_0 = _RAND_752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_1892_1 = _RAND_753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_1892_2 = _RAND_754[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_1892_3 = _RAND_755[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_1902_0 = _RAND_756[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_1902_1 = _RAND_757[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_1902_2 = _RAND_758[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_1902_3 = _RAND_759[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_1912_0 = _RAND_760[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_1912_1 = _RAND_761[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_1912_2 = _RAND_762[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  _T_1912_3 = _RAND_763[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  _T_1922_0 = _RAND_764[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_1922_1 = _RAND_765[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_1922_2 = _RAND_766[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_1922_3 = _RAND_767[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_1932_0 = _RAND_768[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_1932_1 = _RAND_769[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_1932_2 = _RAND_770[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_1932_3 = _RAND_771[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_1942_0 = _RAND_772[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_1942_1 = _RAND_773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_1942_2 = _RAND_774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_1942_3 = _RAND_775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_1952_0 = _RAND_776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_1952_1 = _RAND_777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_1952_2 = _RAND_778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_1952_3 = _RAND_779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_1962_0 = _RAND_780[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_1962_1 = _RAND_781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_1962_2 = _RAND_782[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_1962_3 = _RAND_783[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_1972_0 = _RAND_784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_1972_1 = _RAND_785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_1972_2 = _RAND_786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_1972_3 = _RAND_787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_1982_0 = _RAND_788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_1982_1 = _RAND_789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_1982_2 = _RAND_790[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_1982_3 = _RAND_791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_1992_0 = _RAND_792[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_1992_1 = _RAND_793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_1992_2 = _RAND_794[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_1992_3 = _RAND_795[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_2002_0 = _RAND_796[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_2002_1 = _RAND_797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_2002_2 = _RAND_798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_2002_3 = _RAND_799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_2012_0 = _RAND_800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_2012_1 = _RAND_801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_2012_2 = _RAND_802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_2012_3 = _RAND_803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_2022_0 = _RAND_804[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_2022_1 = _RAND_805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_2022_2 = _RAND_806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_2022_3 = _RAND_807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_2032_0 = _RAND_808[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_2032_1 = _RAND_809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_2032_2 = _RAND_810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_2032_3 = _RAND_811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_2042_0 = _RAND_812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_2042_1 = _RAND_813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_2042_2 = _RAND_814[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_2042_3 = _RAND_815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_2052_0 = _RAND_816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_2052_1 = _RAND_817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_2052_2 = _RAND_818[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_2052_3 = _RAND_819[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_2062_0 = _RAND_820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_2062_1 = _RAND_821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_2062_2 = _RAND_822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_2062_3 = _RAND_823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_2072_0 = _RAND_824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_2072_1 = _RAND_825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_2072_2 = _RAND_826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_2072_3 = _RAND_827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_2082_0 = _RAND_828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_2082_1 = _RAND_829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_2082_2 = _RAND_830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_2082_3 = _RAND_831[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_2092_0 = _RAND_832[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_2092_1 = _RAND_833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_2092_2 = _RAND_834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_2092_3 = _RAND_835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_2102_0 = _RAND_836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_2102_1 = _RAND_837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_2102_2 = _RAND_838[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_2102_3 = _RAND_839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_2112_0 = _RAND_840[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_2112_1 = _RAND_841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_2112_2 = _RAND_842[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_2112_3 = _RAND_843[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_2122_0 = _RAND_844[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_2122_1 = _RAND_845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_2122_2 = _RAND_846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_2122_3 = _RAND_847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_2132_0 = _RAND_848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_2132_1 = _RAND_849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_2132_2 = _RAND_850[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_2132_3 = _RAND_851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_2142_0 = _RAND_852[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_2142_1 = _RAND_853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_2142_2 = _RAND_854[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_2142_3 = _RAND_855[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_2152_0 = _RAND_856[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_2152_1 = _RAND_857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_2152_2 = _RAND_858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_2152_3 = _RAND_859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_2162_0 = _RAND_860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_2162_1 = _RAND_861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_2162_2 = _RAND_862[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_2162_3 = _RAND_863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_2172_0 = _RAND_864[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_2172_1 = _RAND_865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_2172_2 = _RAND_866[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_2172_3 = _RAND_867[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_2182_0 = _RAND_868[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_2182_1 = _RAND_869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_2182_2 = _RAND_870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_2182_3 = _RAND_871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_2192_0 = _RAND_872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_2192_1 = _RAND_873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_2192_2 = _RAND_874[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_2192_3 = _RAND_875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_2202_0 = _RAND_876[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_2202_1 = _RAND_877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_2202_2 = _RAND_878[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_2202_3 = _RAND_879[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_2212_0 = _RAND_880[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_2212_1 = _RAND_881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_2212_2 = _RAND_882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_2212_3 = _RAND_883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_2222_0 = _RAND_884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_2222_1 = _RAND_885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_2222_2 = _RAND_886[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_2222_3 = _RAND_887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_2232_0 = _RAND_888[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_2232_1 = _RAND_889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_2232_2 = _RAND_890[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_2232_3 = _RAND_891[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_2242_0 = _RAND_892[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_2242_1 = _RAND_893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_2242_2 = _RAND_894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_2242_3 = _RAND_895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_2252_0 = _RAND_896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_2252_1 = _RAND_897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_2252_2 = _RAND_898[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_2252_3 = _RAND_899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_2262_0 = _RAND_900[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_2262_1 = _RAND_901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_2262_2 = _RAND_902[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_2262_3 = _RAND_903[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_2272_0 = _RAND_904[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_2272_1 = _RAND_905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_2272_2 = _RAND_906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_2272_3 = _RAND_907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_2282_0 = _RAND_908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_2282_1 = _RAND_909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_2282_2 = _RAND_910[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_2282_3 = _RAND_911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_2292_0 = _RAND_912[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_2292_1 = _RAND_913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_2292_2 = _RAND_914[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_2292_3 = _RAND_915[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_2302_0 = _RAND_916[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_2302_1 = _RAND_917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_2302_2 = _RAND_918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_2302_3 = _RAND_919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_2312_0 = _RAND_920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_2312_1 = _RAND_921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_2312_2 = _RAND_922[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_2312_3 = _RAND_923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_2322_0 = _RAND_924[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_2322_1 = _RAND_925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_2322_2 = _RAND_926[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_2322_3 = _RAND_927[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_2332_0 = _RAND_928[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_2332_1 = _RAND_929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_2332_2 = _RAND_930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_2332_3 = _RAND_931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_2342_0 = _RAND_932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_2342_1 = _RAND_933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_2342_2 = _RAND_934[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_2342_3 = _RAND_935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_2352_0 = _RAND_936[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_2352_1 = _RAND_937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_2352_2 = _RAND_938[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_2352_3 = _RAND_939[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_2362_0 = _RAND_940[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_2362_1 = _RAND_941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_2362_2 = _RAND_942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_2362_3 = _RAND_943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_2372_0 = _RAND_944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_2372_1 = _RAND_945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_2372_2 = _RAND_946[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_2372_3 = _RAND_947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_2382_0 = _RAND_948[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_2382_1 = _RAND_949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_2382_2 = _RAND_950[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_2382_3 = _RAND_951[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_2392_0 = _RAND_952[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_2392_1 = _RAND_953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_2392_2 = _RAND_954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_2392_3 = _RAND_955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_2402_0 = _RAND_956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_2402_1 = _RAND_957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_2402_2 = _RAND_958[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_2402_3 = _RAND_959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_2412_0 = _RAND_960[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_2412_1 = _RAND_961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_2412_2 = _RAND_962[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_2412_3 = _RAND_963[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_2422_0 = _RAND_964[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_2422_1 = _RAND_965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_2422_2 = _RAND_966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_2422_3 = _RAND_967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_2432_0 = _RAND_968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_2432_1 = _RAND_969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_2432_2 = _RAND_970[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_2432_3 = _RAND_971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_2442_0 = _RAND_972[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_2442_1 = _RAND_973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_2442_2 = _RAND_974[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_2442_3 = _RAND_975[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_2452_0 = _RAND_976[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_2452_1 = _RAND_977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_2452_2 = _RAND_978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_2452_3 = _RAND_979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_2462_0 = _RAND_980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_2462_1 = _RAND_981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_2462_2 = _RAND_982[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_2462_3 = _RAND_983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_2472_0 = _RAND_984[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_2472_1 = _RAND_985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_2472_2 = _RAND_986[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_2472_3 = _RAND_987[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_2482_0 = _RAND_988[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_2482_1 = _RAND_989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_2482_2 = _RAND_990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_2482_3 = _RAND_991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_2492_0 = _RAND_992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_2492_1 = _RAND_993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_2492_2 = _RAND_994[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_2492_3 = _RAND_995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_2502_0 = _RAND_996[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_2502_1 = _RAND_997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_2502_2 = _RAND_998[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_2502_3 = _RAND_999[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_2512_0 = _RAND_1000[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_2512_1 = _RAND_1001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_2512_2 = _RAND_1002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_2512_3 = _RAND_1003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_2522_0 = _RAND_1004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_2522_1 = _RAND_1005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_2522_2 = _RAND_1006[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_2522_3 = _RAND_1007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_2532_0 = _RAND_1008[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_2532_1 = _RAND_1009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_2532_2 = _RAND_1010[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_2532_3 = _RAND_1011[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_2542_0 = _RAND_1012[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_2542_1 = _RAND_1013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_2542_2 = _RAND_1014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_2542_3 = _RAND_1015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_2552_0 = _RAND_1016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_2552_1 = _RAND_1017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_2552_2 = _RAND_1018[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_2552_3 = _RAND_1019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_2562_0 = _RAND_1020[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_2562_1 = _RAND_1021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_2562_2 = _RAND_1022[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_2562_3 = _RAND_1023[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_2575_0 = _RAND_1024[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  _T_2575_1 = _RAND_1025[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  _T_2575_2 = _RAND_1026[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  _T_2584_0 = _RAND_1027[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  _T_2584_1 = _RAND_1028[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  _T_2584_2 = _RAND_1029[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  _T_2593_0 = _RAND_1030[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  _T_2593_1 = _RAND_1031[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  _T_2593_2 = _RAND_1032[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  _T_2602_0 = _RAND_1033[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  _T_2602_1 = _RAND_1034[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  _T_2602_2 = _RAND_1035[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  _T_2611_0 = _RAND_1036[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  _T_2611_1 = _RAND_1037[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  _T_2611_2 = _RAND_1038[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  _T_2620_0 = _RAND_1039[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  _T_2620_1 = _RAND_1040[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  _T_2620_2 = _RAND_1041[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  _T_2629_0 = _RAND_1042[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  _T_2629_1 = _RAND_1043[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  _T_2629_2 = _RAND_1044[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  _T_2638_0 = _RAND_1045[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  _T_2638_1 = _RAND_1046[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  _T_2638_2 = _RAND_1047[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  _T_2647_0 = _RAND_1048[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  _T_2647_1 = _RAND_1049[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  _T_2647_2 = _RAND_1050[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  _T_2656_0 = _RAND_1051[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  _T_2656_1 = _RAND_1052[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  _T_2656_2 = _RAND_1053[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  _T_2665_0 = _RAND_1054[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  _T_2665_1 = _RAND_1055[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  _T_2665_2 = _RAND_1056[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  _T_2674_0 = _RAND_1057[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  _T_2674_1 = _RAND_1058[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  _T_2674_2 = _RAND_1059[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  _T_2683_0 = _RAND_1060[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  _T_2683_1 = _RAND_1061[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  _T_2683_2 = _RAND_1062[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  _T_2692_0 = _RAND_1063[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  _T_2692_1 = _RAND_1064[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  _T_2692_2 = _RAND_1065[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  _T_2701_0 = _RAND_1066[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  _T_2701_1 = _RAND_1067[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  _T_2701_2 = _RAND_1068[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  _T_2710_0 = _RAND_1069[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  _T_2710_1 = _RAND_1070[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  _T_2710_2 = _RAND_1071[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  _T_2712_0 = _RAND_1072[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  _T_2712_1 = _RAND_1073[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  _T_2712_2 = _RAND_1074[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  _T_2712_3 = _RAND_1075[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  _T_2712_4 = _RAND_1076[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  _T_2712_5 = _RAND_1077[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  _T_2712_6 = _RAND_1078[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  _T_2712_7 = _RAND_1079[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  _T_2712_8 = _RAND_1080[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  _T_2712_9 = _RAND_1081[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  _T_2712_10 = _RAND_1082[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  _T_2712_11 = _RAND_1083[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  _T_2712_12 = _RAND_1084[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  _T_2712_13 = _RAND_1085[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  _T_2712_14 = _RAND_1086[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  _T_2712_15 = _RAND_1087[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  _T_2712_16 = _RAND_1088[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  _T_2712_17 = _RAND_1089[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  _T_2712_18 = _RAND_1090[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  _T_2712_19 = _RAND_1091[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  _T_2712_20 = _RAND_1092[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  _T_2712_21 = _RAND_1093[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  _T_2712_22 = _RAND_1094[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  _T_2712_23 = _RAND_1095[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  _T_2712_24 = _RAND_1096[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  _T_2712_25 = _RAND_1097[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  _T_2712_26 = _RAND_1098[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  _T_2712_27 = _RAND_1099[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  _T_2712_28 = _RAND_1100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  _T_2712_29 = _RAND_1101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  _T_2712_30 = _RAND_1102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  _T_2712_31 = _RAND_1103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  _T_2712_32 = _RAND_1104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  _T_2712_33 = _RAND_1105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  _T_2712_34 = _RAND_1106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  _T_2712_35 = _RAND_1107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  _T_2712_36 = _RAND_1108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  _T_2712_37 = _RAND_1109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  _T_2712_38 = _RAND_1110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  _T_2712_39 = _RAND_1111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  _T_2712_40 = _RAND_1112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  _T_2712_41 = _RAND_1113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  _T_2712_42 = _RAND_1114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  _T_2712_43 = _RAND_1115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  _T_2712_44 = _RAND_1116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  _T_2712_45 = _RAND_1117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  _T_2712_46 = _RAND_1118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  _T_2712_47 = _RAND_1119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  _T_2712_48 = _RAND_1120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  _T_2712_49 = _RAND_1121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  _T_2712_50 = _RAND_1122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  _T_2712_51 = _RAND_1123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  _T_2712_52 = _RAND_1124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  _T_2712_53 = _RAND_1125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  _T_2712_54 = _RAND_1126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  _T_2712_55 = _RAND_1127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  _T_2712_56 = _RAND_1128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  _T_2712_57 = _RAND_1129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  _T_2712_58 = _RAND_1130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  _T_2712_59 = _RAND_1131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  _T_2712_60 = _RAND_1132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  _T_2712_61 = _RAND_1133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  _T_2712_62 = _RAND_1134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  _T_2712_63 = _RAND_1135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  _T_2712_64 = _RAND_1136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  _T_2712_65 = _RAND_1137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  _T_2712_66 = _RAND_1138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  _T_2712_67 = _RAND_1139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  _T_2712_68 = _RAND_1140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  _T_2712_69 = _RAND_1141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  _T_2712_70 = _RAND_1142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  _T_2712_71 = _RAND_1143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  _T_2712_72 = _RAND_1144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  _T_2712_73 = _RAND_1145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  _T_2712_74 = _RAND_1146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  _T_2712_75 = _RAND_1147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  _T_2712_76 = _RAND_1148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  _T_2712_77 = _RAND_1149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  _T_2712_78 = _RAND_1150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  _T_2712_79 = _RAND_1151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  _T_2712_80 = _RAND_1152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  _T_2712_81 = _RAND_1153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  _T_2712_82 = _RAND_1154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  _T_2712_83 = _RAND_1155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  _T_2712_84 = _RAND_1156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  _T_2712_85 = _RAND_1157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  _T_2712_86 = _RAND_1158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  _T_2712_87 = _RAND_1159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  _T_2712_88 = _RAND_1160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  _T_2712_89 = _RAND_1161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  _T_2712_90 = _RAND_1162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  _T_2712_91 = _RAND_1163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  _T_2712_92 = _RAND_1164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  _T_2712_93 = _RAND_1165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  _T_2712_94 = _RAND_1166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  _T_2712_95 = _RAND_1167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  _T_2712_96 = _RAND_1168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  _T_2712_97 = _RAND_1169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  _T_2712_98 = _RAND_1170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  _T_2712_99 = _RAND_1171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  _T_2712_100 = _RAND_1172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  _T_2712_101 = _RAND_1173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  _T_2712_102 = _RAND_1174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  _T_2712_103 = _RAND_1175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  _T_2712_104 = _RAND_1176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  _T_2712_105 = _RAND_1177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  _T_2712_106 = _RAND_1178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  _T_2712_107 = _RAND_1179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  _T_2712_108 = _RAND_1180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  _T_2712_109 = _RAND_1181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  _T_2712_110 = _RAND_1182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  _T_2712_111 = _RAND_1183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  _T_2712_112 = _RAND_1184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  _T_2712_113 = _RAND_1185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  _T_2712_114 = _RAND_1186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  _T_2712_115 = _RAND_1187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  _T_2712_116 = _RAND_1188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  _T_2712_117 = _RAND_1189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  _T_2712_118 = _RAND_1190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  _T_2712_119 = _RAND_1191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  _T_2712_120 = _RAND_1192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  _T_2712_121 = _RAND_1193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  _T_2712_122 = _RAND_1194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  _T_2712_123 = _RAND_1195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  _T_2712_124 = _RAND_1196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  _T_2712_125 = _RAND_1197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  _T_2712_126 = _RAND_1198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  _T_2712_127 = _RAND_1199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  _T_2712_128 = _RAND_1200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  _T_2712_129 = _RAND_1201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  _T_2712_130 = _RAND_1202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  _T_2712_131 = _RAND_1203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  _T_2712_132 = _RAND_1204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  _T_2712_133 = _RAND_1205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  _T_2712_134 = _RAND_1206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  _T_2712_135 = _RAND_1207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  _T_2712_136 = _RAND_1208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  _T_2712_137 = _RAND_1209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  _T_2712_138 = _RAND_1210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  _T_2712_139 = _RAND_1211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  _T_2712_140 = _RAND_1212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  _T_2712_141 = _RAND_1213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  _T_2712_142 = _RAND_1214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  _T_2712_143 = _RAND_1215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  _T_2712_144 = _RAND_1216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  _T_2712_145 = _RAND_1217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  _T_2712_146 = _RAND_1218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  _T_2712_147 = _RAND_1219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  _T_2712_148 = _RAND_1220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  _T_2712_149 = _RAND_1221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  _T_2712_150 = _RAND_1222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  _T_2712_151 = _RAND_1223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  _T_2712_152 = _RAND_1224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  _T_2712_153 = _RAND_1225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  _T_2712_154 = _RAND_1226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  _T_2712_155 = _RAND_1227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  _T_2712_156 = _RAND_1228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  _T_2712_157 = _RAND_1229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  _T_2712_158 = _RAND_1230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  _T_2712_159 = _RAND_1231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  _T_2712_160 = _RAND_1232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  _T_2712_161 = _RAND_1233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  _T_2712_162 = _RAND_1234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  _T_2712_163 = _RAND_1235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  _T_2712_164 = _RAND_1236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  _T_2712_165 = _RAND_1237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  _T_2712_166 = _RAND_1238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  _T_2712_167 = _RAND_1239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  _T_2712_168 = _RAND_1240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  _T_2712_169 = _RAND_1241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  _T_2712_170 = _RAND_1242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  _T_2712_171 = _RAND_1243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  _T_2712_172 = _RAND_1244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  _T_2712_173 = _RAND_1245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  _T_2712_174 = _RAND_1246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  _T_2712_175 = _RAND_1247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  _T_2712_176 = _RAND_1248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  _T_2712_177 = _RAND_1249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  _T_2712_178 = _RAND_1250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  _T_2712_179 = _RAND_1251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_12_0 <= 1'h0;
    end else begin
      _T_12_0 <= _T_5;
    end
    if (reset) begin
      _T_12_1 <= 1'h0;
    end else begin
      _T_12_1 <= _T_12_0;
    end
    if (reset) begin
      _T_12_2 <= 1'h0;
    end else begin
      _T_12_2 <= _T_12_1;
    end
    if (reset) begin
      _T_12_3 <= 1'h0;
    end else begin
      _T_12_3 <= _T_12_2;
    end
    if (reset) begin
      _T_22_0 <= 1'h0;
    end else begin
      _T_22_0 <= _T_15;
    end
    if (reset) begin
      _T_22_1 <= 1'h0;
    end else begin
      _T_22_1 <= _T_22_0;
    end
    if (reset) begin
      _T_22_2 <= 1'h0;
    end else begin
      _T_22_2 <= _T_22_1;
    end
    if (reset) begin
      _T_22_3 <= 1'h0;
    end else begin
      _T_22_3 <= _T_22_2;
    end
    if (reset) begin
      _T_32_0 <= 1'h0;
    end else begin
      _T_32_0 <= _T_25;
    end
    if (reset) begin
      _T_32_1 <= 1'h0;
    end else begin
      _T_32_1 <= _T_32_0;
    end
    if (reset) begin
      _T_32_2 <= 1'h0;
    end else begin
      _T_32_2 <= _T_32_1;
    end
    if (reset) begin
      _T_32_3 <= 1'h0;
    end else begin
      _T_32_3 <= _T_32_2;
    end
    if (reset) begin
      _T_42_0 <= 1'h0;
    end else begin
      _T_42_0 <= _T_35;
    end
    if (reset) begin
      _T_42_1 <= 1'h0;
    end else begin
      _T_42_1 <= _T_42_0;
    end
    if (reset) begin
      _T_42_2 <= 1'h0;
    end else begin
      _T_42_2 <= _T_42_1;
    end
    if (reset) begin
      _T_42_3 <= 1'h0;
    end else begin
      _T_42_3 <= _T_42_2;
    end
    if (reset) begin
      _T_52_0 <= 1'h0;
    end else begin
      _T_52_0 <= _T_45;
    end
    if (reset) begin
      _T_52_1 <= 1'h0;
    end else begin
      _T_52_1 <= _T_52_0;
    end
    if (reset) begin
      _T_52_2 <= 1'h0;
    end else begin
      _T_52_2 <= _T_52_1;
    end
    if (reset) begin
      _T_52_3 <= 1'h0;
    end else begin
      _T_52_3 <= _T_52_2;
    end
    if (reset) begin
      _T_62_0 <= 1'h0;
    end else begin
      _T_62_0 <= _T_55;
    end
    if (reset) begin
      _T_62_1 <= 1'h0;
    end else begin
      _T_62_1 <= _T_62_0;
    end
    if (reset) begin
      _T_62_2 <= 1'h0;
    end else begin
      _T_62_2 <= _T_62_1;
    end
    if (reset) begin
      _T_62_3 <= 1'h0;
    end else begin
      _T_62_3 <= _T_62_2;
    end
    if (reset) begin
      _T_72_0 <= 1'h0;
    end else begin
      _T_72_0 <= _T_65;
    end
    if (reset) begin
      _T_72_1 <= 1'h0;
    end else begin
      _T_72_1 <= _T_72_0;
    end
    if (reset) begin
      _T_72_2 <= 1'h0;
    end else begin
      _T_72_2 <= _T_72_1;
    end
    if (reset) begin
      _T_72_3 <= 1'h0;
    end else begin
      _T_72_3 <= _T_72_2;
    end
    if (reset) begin
      _T_82_0 <= 1'h0;
    end else begin
      _T_82_0 <= _T_75;
    end
    if (reset) begin
      _T_82_1 <= 1'h0;
    end else begin
      _T_82_1 <= _T_82_0;
    end
    if (reset) begin
      _T_82_2 <= 1'h0;
    end else begin
      _T_82_2 <= _T_82_1;
    end
    if (reset) begin
      _T_82_3 <= 1'h0;
    end else begin
      _T_82_3 <= _T_82_2;
    end
    if (reset) begin
      _T_92_0 <= 1'h0;
    end else begin
      _T_92_0 <= _T_85;
    end
    if (reset) begin
      _T_92_1 <= 1'h0;
    end else begin
      _T_92_1 <= _T_92_0;
    end
    if (reset) begin
      _T_92_2 <= 1'h0;
    end else begin
      _T_92_2 <= _T_92_1;
    end
    if (reset) begin
      _T_92_3 <= 1'h0;
    end else begin
      _T_92_3 <= _T_92_2;
    end
    if (reset) begin
      _T_102_0 <= 1'h0;
    end else begin
      _T_102_0 <= _T_95;
    end
    if (reset) begin
      _T_102_1 <= 1'h0;
    end else begin
      _T_102_1 <= _T_102_0;
    end
    if (reset) begin
      _T_102_2 <= 1'h0;
    end else begin
      _T_102_2 <= _T_102_1;
    end
    if (reset) begin
      _T_102_3 <= 1'h0;
    end else begin
      _T_102_3 <= _T_102_2;
    end
    if (reset) begin
      _T_112_0 <= 1'h0;
    end else begin
      _T_112_0 <= _T_105;
    end
    if (reset) begin
      _T_112_1 <= 1'h0;
    end else begin
      _T_112_1 <= _T_112_0;
    end
    if (reset) begin
      _T_112_2 <= 1'h0;
    end else begin
      _T_112_2 <= _T_112_1;
    end
    if (reset) begin
      _T_112_3 <= 1'h0;
    end else begin
      _T_112_3 <= _T_112_2;
    end
    if (reset) begin
      _T_122_0 <= 1'h0;
    end else begin
      _T_122_0 <= _T_115;
    end
    if (reset) begin
      _T_122_1 <= 1'h0;
    end else begin
      _T_122_1 <= _T_122_0;
    end
    if (reset) begin
      _T_122_2 <= 1'h0;
    end else begin
      _T_122_2 <= _T_122_1;
    end
    if (reset) begin
      _T_122_3 <= 1'h0;
    end else begin
      _T_122_3 <= _T_122_2;
    end
    if (reset) begin
      _T_132_0 <= 1'h0;
    end else begin
      _T_132_0 <= _T_125;
    end
    if (reset) begin
      _T_132_1 <= 1'h0;
    end else begin
      _T_132_1 <= _T_132_0;
    end
    if (reset) begin
      _T_132_2 <= 1'h0;
    end else begin
      _T_132_2 <= _T_132_1;
    end
    if (reset) begin
      _T_132_3 <= 1'h0;
    end else begin
      _T_132_3 <= _T_132_2;
    end
    if (reset) begin
      _T_142_0 <= 1'h0;
    end else begin
      _T_142_0 <= _T_135;
    end
    if (reset) begin
      _T_142_1 <= 1'h0;
    end else begin
      _T_142_1 <= _T_142_0;
    end
    if (reset) begin
      _T_142_2 <= 1'h0;
    end else begin
      _T_142_2 <= _T_142_1;
    end
    if (reset) begin
      _T_142_3 <= 1'h0;
    end else begin
      _T_142_3 <= _T_142_2;
    end
    if (reset) begin
      _T_152_0 <= 1'h0;
    end else begin
      _T_152_0 <= _T_145;
    end
    if (reset) begin
      _T_152_1 <= 1'h0;
    end else begin
      _T_152_1 <= _T_152_0;
    end
    if (reset) begin
      _T_152_2 <= 1'h0;
    end else begin
      _T_152_2 <= _T_152_1;
    end
    if (reset) begin
      _T_152_3 <= 1'h0;
    end else begin
      _T_152_3 <= _T_152_2;
    end
    if (reset) begin
      _T_162_0 <= 1'h0;
    end else begin
      _T_162_0 <= _T_155;
    end
    if (reset) begin
      _T_162_1 <= 1'h0;
    end else begin
      _T_162_1 <= _T_162_0;
    end
    if (reset) begin
      _T_162_2 <= 1'h0;
    end else begin
      _T_162_2 <= _T_162_1;
    end
    if (reset) begin
      _T_162_3 <= 1'h0;
    end else begin
      _T_162_3 <= _T_162_2;
    end
    if (reset) begin
      _T_172_0 <= 1'h0;
    end else begin
      _T_172_0 <= _T_15;
    end
    if (reset) begin
      _T_172_1 <= 1'h0;
    end else begin
      _T_172_1 <= _T_172_0;
    end
    if (reset) begin
      _T_172_2 <= 1'h0;
    end else begin
      _T_172_2 <= _T_172_1;
    end
    if (reset) begin
      _T_172_3 <= 1'h0;
    end else begin
      _T_172_3 <= _T_172_2;
    end
    if (reset) begin
      _T_182_0 <= 1'h0;
    end else begin
      _T_182_0 <= _T_25;
    end
    if (reset) begin
      _T_182_1 <= 1'h0;
    end else begin
      _T_182_1 <= _T_182_0;
    end
    if (reset) begin
      _T_182_2 <= 1'h0;
    end else begin
      _T_182_2 <= _T_182_1;
    end
    if (reset) begin
      _T_182_3 <= 1'h0;
    end else begin
      _T_182_3 <= _T_182_2;
    end
    if (reset) begin
      _T_192_0 <= 1'h0;
    end else begin
      _T_192_0 <= _T_35;
    end
    if (reset) begin
      _T_192_1 <= 1'h0;
    end else begin
      _T_192_1 <= _T_192_0;
    end
    if (reset) begin
      _T_192_2 <= 1'h0;
    end else begin
      _T_192_2 <= _T_192_1;
    end
    if (reset) begin
      _T_192_3 <= 1'h0;
    end else begin
      _T_192_3 <= _T_192_2;
    end
    if (reset) begin
      _T_202_0 <= 1'h0;
    end else begin
      _T_202_0 <= _T_45;
    end
    if (reset) begin
      _T_202_1 <= 1'h0;
    end else begin
      _T_202_1 <= _T_202_0;
    end
    if (reset) begin
      _T_202_2 <= 1'h0;
    end else begin
      _T_202_2 <= _T_202_1;
    end
    if (reset) begin
      _T_202_3 <= 1'h0;
    end else begin
      _T_202_3 <= _T_202_2;
    end
    if (reset) begin
      _T_212_0 <= 1'h0;
    end else begin
      _T_212_0 <= _T_55;
    end
    if (reset) begin
      _T_212_1 <= 1'h0;
    end else begin
      _T_212_1 <= _T_212_0;
    end
    if (reset) begin
      _T_212_2 <= 1'h0;
    end else begin
      _T_212_2 <= _T_212_1;
    end
    if (reset) begin
      _T_212_3 <= 1'h0;
    end else begin
      _T_212_3 <= _T_212_2;
    end
    if (reset) begin
      _T_222_0 <= 1'h0;
    end else begin
      _T_222_0 <= _T_65;
    end
    if (reset) begin
      _T_222_1 <= 1'h0;
    end else begin
      _T_222_1 <= _T_222_0;
    end
    if (reset) begin
      _T_222_2 <= 1'h0;
    end else begin
      _T_222_2 <= _T_222_1;
    end
    if (reset) begin
      _T_222_3 <= 1'h0;
    end else begin
      _T_222_3 <= _T_222_2;
    end
    if (reset) begin
      _T_232_0 <= 1'h0;
    end else begin
      _T_232_0 <= _T_75;
    end
    if (reset) begin
      _T_232_1 <= 1'h0;
    end else begin
      _T_232_1 <= _T_232_0;
    end
    if (reset) begin
      _T_232_2 <= 1'h0;
    end else begin
      _T_232_2 <= _T_232_1;
    end
    if (reset) begin
      _T_232_3 <= 1'h0;
    end else begin
      _T_232_3 <= _T_232_2;
    end
    if (reset) begin
      _T_242_0 <= 1'h0;
    end else begin
      _T_242_0 <= _T_85;
    end
    if (reset) begin
      _T_242_1 <= 1'h0;
    end else begin
      _T_242_1 <= _T_242_0;
    end
    if (reset) begin
      _T_242_2 <= 1'h0;
    end else begin
      _T_242_2 <= _T_242_1;
    end
    if (reset) begin
      _T_242_3 <= 1'h0;
    end else begin
      _T_242_3 <= _T_242_2;
    end
    if (reset) begin
      _T_252_0 <= 1'h0;
    end else begin
      _T_252_0 <= _T_95;
    end
    if (reset) begin
      _T_252_1 <= 1'h0;
    end else begin
      _T_252_1 <= _T_252_0;
    end
    if (reset) begin
      _T_252_2 <= 1'h0;
    end else begin
      _T_252_2 <= _T_252_1;
    end
    if (reset) begin
      _T_252_3 <= 1'h0;
    end else begin
      _T_252_3 <= _T_252_2;
    end
    if (reset) begin
      _T_262_0 <= 1'h0;
    end else begin
      _T_262_0 <= _T_105;
    end
    if (reset) begin
      _T_262_1 <= 1'h0;
    end else begin
      _T_262_1 <= _T_262_0;
    end
    if (reset) begin
      _T_262_2 <= 1'h0;
    end else begin
      _T_262_2 <= _T_262_1;
    end
    if (reset) begin
      _T_262_3 <= 1'h0;
    end else begin
      _T_262_3 <= _T_262_2;
    end
    if (reset) begin
      _T_272_0 <= 1'h0;
    end else begin
      _T_272_0 <= _T_115;
    end
    if (reset) begin
      _T_272_1 <= 1'h0;
    end else begin
      _T_272_1 <= _T_272_0;
    end
    if (reset) begin
      _T_272_2 <= 1'h0;
    end else begin
      _T_272_2 <= _T_272_1;
    end
    if (reset) begin
      _T_272_3 <= 1'h0;
    end else begin
      _T_272_3 <= _T_272_2;
    end
    if (reset) begin
      _T_282_0 <= 1'h0;
    end else begin
      _T_282_0 <= _T_125;
    end
    if (reset) begin
      _T_282_1 <= 1'h0;
    end else begin
      _T_282_1 <= _T_282_0;
    end
    if (reset) begin
      _T_282_2 <= 1'h0;
    end else begin
      _T_282_2 <= _T_282_1;
    end
    if (reset) begin
      _T_282_3 <= 1'h0;
    end else begin
      _T_282_3 <= _T_282_2;
    end
    if (reset) begin
      _T_292_0 <= 1'h0;
    end else begin
      _T_292_0 <= _T_135;
    end
    if (reset) begin
      _T_292_1 <= 1'h0;
    end else begin
      _T_292_1 <= _T_292_0;
    end
    if (reset) begin
      _T_292_2 <= 1'h0;
    end else begin
      _T_292_2 <= _T_292_1;
    end
    if (reset) begin
      _T_292_3 <= 1'h0;
    end else begin
      _T_292_3 <= _T_292_2;
    end
    if (reset) begin
      _T_302_0 <= 1'h0;
    end else begin
      _T_302_0 <= _T_145;
    end
    if (reset) begin
      _T_302_1 <= 1'h0;
    end else begin
      _T_302_1 <= _T_302_0;
    end
    if (reset) begin
      _T_302_2 <= 1'h0;
    end else begin
      _T_302_2 <= _T_302_1;
    end
    if (reset) begin
      _T_302_3 <= 1'h0;
    end else begin
      _T_302_3 <= _T_302_2;
    end
    if (reset) begin
      _T_312_0 <= 1'h0;
    end else begin
      _T_312_0 <= _T_155;
    end
    if (reset) begin
      _T_312_1 <= 1'h0;
    end else begin
      _T_312_1 <= _T_312_0;
    end
    if (reset) begin
      _T_312_2 <= 1'h0;
    end else begin
      _T_312_2 <= _T_312_1;
    end
    if (reset) begin
      _T_312_3 <= 1'h0;
    end else begin
      _T_312_3 <= _T_312_2;
    end
    if (reset) begin
      _T_322_0 <= 1'h0;
    end else begin
      _T_322_0 <= _T_315;
    end
    if (reset) begin
      _T_322_1 <= 1'h0;
    end else begin
      _T_322_1 <= _T_322_0;
    end
    if (reset) begin
      _T_322_2 <= 1'h0;
    end else begin
      _T_322_2 <= _T_322_1;
    end
    if (reset) begin
      _T_322_3 <= 1'h0;
    end else begin
      _T_322_3 <= _T_322_2;
    end
    if (reset) begin
      _T_332_0 <= 1'h0;
    end else begin
      _T_332_0 <= _T_25;
    end
    if (reset) begin
      _T_332_1 <= 1'h0;
    end else begin
      _T_332_1 <= _T_332_0;
    end
    if (reset) begin
      _T_332_2 <= 1'h0;
    end else begin
      _T_332_2 <= _T_332_1;
    end
    if (reset) begin
      _T_332_3 <= 1'h0;
    end else begin
      _T_332_3 <= _T_332_2;
    end
    if (reset) begin
      _T_342_0 <= 1'h0;
    end else begin
      _T_342_0 <= _T_35;
    end
    if (reset) begin
      _T_342_1 <= 1'h0;
    end else begin
      _T_342_1 <= _T_342_0;
    end
    if (reset) begin
      _T_342_2 <= 1'h0;
    end else begin
      _T_342_2 <= _T_342_1;
    end
    if (reset) begin
      _T_342_3 <= 1'h0;
    end else begin
      _T_342_3 <= _T_342_2;
    end
    if (reset) begin
      _T_352_0 <= 1'h0;
    end else begin
      _T_352_0 <= _T_45;
    end
    if (reset) begin
      _T_352_1 <= 1'h0;
    end else begin
      _T_352_1 <= _T_352_0;
    end
    if (reset) begin
      _T_352_2 <= 1'h0;
    end else begin
      _T_352_2 <= _T_352_1;
    end
    if (reset) begin
      _T_352_3 <= 1'h0;
    end else begin
      _T_352_3 <= _T_352_2;
    end
    if (reset) begin
      _T_362_0 <= 1'h0;
    end else begin
      _T_362_0 <= _T_55;
    end
    if (reset) begin
      _T_362_1 <= 1'h0;
    end else begin
      _T_362_1 <= _T_362_0;
    end
    if (reset) begin
      _T_362_2 <= 1'h0;
    end else begin
      _T_362_2 <= _T_362_1;
    end
    if (reset) begin
      _T_362_3 <= 1'h0;
    end else begin
      _T_362_3 <= _T_362_2;
    end
    if (reset) begin
      _T_372_0 <= 1'h0;
    end else begin
      _T_372_0 <= _T_65;
    end
    if (reset) begin
      _T_372_1 <= 1'h0;
    end else begin
      _T_372_1 <= _T_372_0;
    end
    if (reset) begin
      _T_372_2 <= 1'h0;
    end else begin
      _T_372_2 <= _T_372_1;
    end
    if (reset) begin
      _T_372_3 <= 1'h0;
    end else begin
      _T_372_3 <= _T_372_2;
    end
    if (reset) begin
      _T_382_0 <= 1'h0;
    end else begin
      _T_382_0 <= _T_75;
    end
    if (reset) begin
      _T_382_1 <= 1'h0;
    end else begin
      _T_382_1 <= _T_382_0;
    end
    if (reset) begin
      _T_382_2 <= 1'h0;
    end else begin
      _T_382_2 <= _T_382_1;
    end
    if (reset) begin
      _T_382_3 <= 1'h0;
    end else begin
      _T_382_3 <= _T_382_2;
    end
    if (reset) begin
      _T_392_0 <= 1'h0;
    end else begin
      _T_392_0 <= _T_85;
    end
    if (reset) begin
      _T_392_1 <= 1'h0;
    end else begin
      _T_392_1 <= _T_392_0;
    end
    if (reset) begin
      _T_392_2 <= 1'h0;
    end else begin
      _T_392_2 <= _T_392_1;
    end
    if (reset) begin
      _T_392_3 <= 1'h0;
    end else begin
      _T_392_3 <= _T_392_2;
    end
    if (reset) begin
      _T_402_0 <= 1'h0;
    end else begin
      _T_402_0 <= _T_95;
    end
    if (reset) begin
      _T_402_1 <= 1'h0;
    end else begin
      _T_402_1 <= _T_402_0;
    end
    if (reset) begin
      _T_402_2 <= 1'h0;
    end else begin
      _T_402_2 <= _T_402_1;
    end
    if (reset) begin
      _T_402_3 <= 1'h0;
    end else begin
      _T_402_3 <= _T_402_2;
    end
    if (reset) begin
      _T_412_0 <= 1'h0;
    end else begin
      _T_412_0 <= _T_105;
    end
    if (reset) begin
      _T_412_1 <= 1'h0;
    end else begin
      _T_412_1 <= _T_412_0;
    end
    if (reset) begin
      _T_412_2 <= 1'h0;
    end else begin
      _T_412_2 <= _T_412_1;
    end
    if (reset) begin
      _T_412_3 <= 1'h0;
    end else begin
      _T_412_3 <= _T_412_2;
    end
    if (reset) begin
      _T_422_0 <= 1'h0;
    end else begin
      _T_422_0 <= _T_115;
    end
    if (reset) begin
      _T_422_1 <= 1'h0;
    end else begin
      _T_422_1 <= _T_422_0;
    end
    if (reset) begin
      _T_422_2 <= 1'h0;
    end else begin
      _T_422_2 <= _T_422_1;
    end
    if (reset) begin
      _T_422_3 <= 1'h0;
    end else begin
      _T_422_3 <= _T_422_2;
    end
    if (reset) begin
      _T_432_0 <= 1'h0;
    end else begin
      _T_432_0 <= _T_125;
    end
    if (reset) begin
      _T_432_1 <= 1'h0;
    end else begin
      _T_432_1 <= _T_432_0;
    end
    if (reset) begin
      _T_432_2 <= 1'h0;
    end else begin
      _T_432_2 <= _T_432_1;
    end
    if (reset) begin
      _T_432_3 <= 1'h0;
    end else begin
      _T_432_3 <= _T_432_2;
    end
    if (reset) begin
      _T_442_0 <= 1'h0;
    end else begin
      _T_442_0 <= _T_135;
    end
    if (reset) begin
      _T_442_1 <= 1'h0;
    end else begin
      _T_442_1 <= _T_442_0;
    end
    if (reset) begin
      _T_442_2 <= 1'h0;
    end else begin
      _T_442_2 <= _T_442_1;
    end
    if (reset) begin
      _T_442_3 <= 1'h0;
    end else begin
      _T_442_3 <= _T_442_2;
    end
    if (reset) begin
      _T_452_0 <= 1'h0;
    end else begin
      _T_452_0 <= _T_145;
    end
    if (reset) begin
      _T_452_1 <= 1'h0;
    end else begin
      _T_452_1 <= _T_452_0;
    end
    if (reset) begin
      _T_452_2 <= 1'h0;
    end else begin
      _T_452_2 <= _T_452_1;
    end
    if (reset) begin
      _T_452_3 <= 1'h0;
    end else begin
      _T_452_3 <= _T_452_2;
    end
    if (reset) begin
      _T_462_0 <= 1'h0;
    end else begin
      _T_462_0 <= _T_155;
    end
    if (reset) begin
      _T_462_1 <= 1'h0;
    end else begin
      _T_462_1 <= _T_462_0;
    end
    if (reset) begin
      _T_462_2 <= 1'h0;
    end else begin
      _T_462_2 <= _T_462_1;
    end
    if (reset) begin
      _T_462_3 <= 1'h0;
    end else begin
      _T_462_3 <= _T_462_2;
    end
    if (reset) begin
      _T_472_0 <= 1'h0;
    end else begin
      _T_472_0 <= _T_315;
    end
    if (reset) begin
      _T_472_1 <= 1'h0;
    end else begin
      _T_472_1 <= _T_472_0;
    end
    if (reset) begin
      _T_472_2 <= 1'h0;
    end else begin
      _T_472_2 <= _T_472_1;
    end
    if (reset) begin
      _T_472_3 <= 1'h0;
    end else begin
      _T_472_3 <= _T_472_2;
    end
    if (reset) begin
      _T_482_0 <= 1'h0;
    end else begin
      _T_482_0 <= _T_475;
    end
    if (reset) begin
      _T_482_1 <= 1'h0;
    end else begin
      _T_482_1 <= _T_482_0;
    end
    if (reset) begin
      _T_482_2 <= 1'h0;
    end else begin
      _T_482_2 <= _T_482_1;
    end
    if (reset) begin
      _T_482_3 <= 1'h0;
    end else begin
      _T_482_3 <= _T_482_2;
    end
    if (reset) begin
      _T_492_0 <= 1'h0;
    end else begin
      _T_492_0 <= _T_35;
    end
    if (reset) begin
      _T_492_1 <= 1'h0;
    end else begin
      _T_492_1 <= _T_492_0;
    end
    if (reset) begin
      _T_492_2 <= 1'h0;
    end else begin
      _T_492_2 <= _T_492_1;
    end
    if (reset) begin
      _T_492_3 <= 1'h0;
    end else begin
      _T_492_3 <= _T_492_2;
    end
    if (reset) begin
      _T_502_0 <= 1'h0;
    end else begin
      _T_502_0 <= _T_45;
    end
    if (reset) begin
      _T_502_1 <= 1'h0;
    end else begin
      _T_502_1 <= _T_502_0;
    end
    if (reset) begin
      _T_502_2 <= 1'h0;
    end else begin
      _T_502_2 <= _T_502_1;
    end
    if (reset) begin
      _T_502_3 <= 1'h0;
    end else begin
      _T_502_3 <= _T_502_2;
    end
    if (reset) begin
      _T_512_0 <= 1'h0;
    end else begin
      _T_512_0 <= _T_55;
    end
    if (reset) begin
      _T_512_1 <= 1'h0;
    end else begin
      _T_512_1 <= _T_512_0;
    end
    if (reset) begin
      _T_512_2 <= 1'h0;
    end else begin
      _T_512_2 <= _T_512_1;
    end
    if (reset) begin
      _T_512_3 <= 1'h0;
    end else begin
      _T_512_3 <= _T_512_2;
    end
    if (reset) begin
      _T_522_0 <= 1'h0;
    end else begin
      _T_522_0 <= _T_65;
    end
    if (reset) begin
      _T_522_1 <= 1'h0;
    end else begin
      _T_522_1 <= _T_522_0;
    end
    if (reset) begin
      _T_522_2 <= 1'h0;
    end else begin
      _T_522_2 <= _T_522_1;
    end
    if (reset) begin
      _T_522_3 <= 1'h0;
    end else begin
      _T_522_3 <= _T_522_2;
    end
    if (reset) begin
      _T_532_0 <= 1'h0;
    end else begin
      _T_532_0 <= _T_75;
    end
    if (reset) begin
      _T_532_1 <= 1'h0;
    end else begin
      _T_532_1 <= _T_532_0;
    end
    if (reset) begin
      _T_532_2 <= 1'h0;
    end else begin
      _T_532_2 <= _T_532_1;
    end
    if (reset) begin
      _T_532_3 <= 1'h0;
    end else begin
      _T_532_3 <= _T_532_2;
    end
    if (reset) begin
      _T_542_0 <= 1'h0;
    end else begin
      _T_542_0 <= _T_85;
    end
    if (reset) begin
      _T_542_1 <= 1'h0;
    end else begin
      _T_542_1 <= _T_542_0;
    end
    if (reset) begin
      _T_542_2 <= 1'h0;
    end else begin
      _T_542_2 <= _T_542_1;
    end
    if (reset) begin
      _T_542_3 <= 1'h0;
    end else begin
      _T_542_3 <= _T_542_2;
    end
    if (reset) begin
      _T_552_0 <= 1'h0;
    end else begin
      _T_552_0 <= _T_95;
    end
    if (reset) begin
      _T_552_1 <= 1'h0;
    end else begin
      _T_552_1 <= _T_552_0;
    end
    if (reset) begin
      _T_552_2 <= 1'h0;
    end else begin
      _T_552_2 <= _T_552_1;
    end
    if (reset) begin
      _T_552_3 <= 1'h0;
    end else begin
      _T_552_3 <= _T_552_2;
    end
    if (reset) begin
      _T_562_0 <= 1'h0;
    end else begin
      _T_562_0 <= _T_105;
    end
    if (reset) begin
      _T_562_1 <= 1'h0;
    end else begin
      _T_562_1 <= _T_562_0;
    end
    if (reset) begin
      _T_562_2 <= 1'h0;
    end else begin
      _T_562_2 <= _T_562_1;
    end
    if (reset) begin
      _T_562_3 <= 1'h0;
    end else begin
      _T_562_3 <= _T_562_2;
    end
    if (reset) begin
      _T_572_0 <= 1'h0;
    end else begin
      _T_572_0 <= _T_115;
    end
    if (reset) begin
      _T_572_1 <= 1'h0;
    end else begin
      _T_572_1 <= _T_572_0;
    end
    if (reset) begin
      _T_572_2 <= 1'h0;
    end else begin
      _T_572_2 <= _T_572_1;
    end
    if (reset) begin
      _T_572_3 <= 1'h0;
    end else begin
      _T_572_3 <= _T_572_2;
    end
    if (reset) begin
      _T_582_0 <= 1'h0;
    end else begin
      _T_582_0 <= _T_125;
    end
    if (reset) begin
      _T_582_1 <= 1'h0;
    end else begin
      _T_582_1 <= _T_582_0;
    end
    if (reset) begin
      _T_582_2 <= 1'h0;
    end else begin
      _T_582_2 <= _T_582_1;
    end
    if (reset) begin
      _T_582_3 <= 1'h0;
    end else begin
      _T_582_3 <= _T_582_2;
    end
    if (reset) begin
      _T_592_0 <= 1'h0;
    end else begin
      _T_592_0 <= _T_135;
    end
    if (reset) begin
      _T_592_1 <= 1'h0;
    end else begin
      _T_592_1 <= _T_592_0;
    end
    if (reset) begin
      _T_592_2 <= 1'h0;
    end else begin
      _T_592_2 <= _T_592_1;
    end
    if (reset) begin
      _T_592_3 <= 1'h0;
    end else begin
      _T_592_3 <= _T_592_2;
    end
    if (reset) begin
      _T_602_0 <= 1'h0;
    end else begin
      _T_602_0 <= _T_145;
    end
    if (reset) begin
      _T_602_1 <= 1'h0;
    end else begin
      _T_602_1 <= _T_602_0;
    end
    if (reset) begin
      _T_602_2 <= 1'h0;
    end else begin
      _T_602_2 <= _T_602_1;
    end
    if (reset) begin
      _T_602_3 <= 1'h0;
    end else begin
      _T_602_3 <= _T_602_2;
    end
    if (reset) begin
      _T_612_0 <= 1'h0;
    end else begin
      _T_612_0 <= _T_155;
    end
    if (reset) begin
      _T_612_1 <= 1'h0;
    end else begin
      _T_612_1 <= _T_612_0;
    end
    if (reset) begin
      _T_612_2 <= 1'h0;
    end else begin
      _T_612_2 <= _T_612_1;
    end
    if (reset) begin
      _T_612_3 <= 1'h0;
    end else begin
      _T_612_3 <= _T_612_2;
    end
    if (reset) begin
      _T_622_0 <= 1'h0;
    end else begin
      _T_622_0 <= _T_315;
    end
    if (reset) begin
      _T_622_1 <= 1'h0;
    end else begin
      _T_622_1 <= _T_622_0;
    end
    if (reset) begin
      _T_622_2 <= 1'h0;
    end else begin
      _T_622_2 <= _T_622_1;
    end
    if (reset) begin
      _T_622_3 <= 1'h0;
    end else begin
      _T_622_3 <= _T_622_2;
    end
    if (reset) begin
      _T_632_0 <= 1'h0;
    end else begin
      _T_632_0 <= _T_475;
    end
    if (reset) begin
      _T_632_1 <= 1'h0;
    end else begin
      _T_632_1 <= _T_632_0;
    end
    if (reset) begin
      _T_632_2 <= 1'h0;
    end else begin
      _T_632_2 <= _T_632_1;
    end
    if (reset) begin
      _T_632_3 <= 1'h0;
    end else begin
      _T_632_3 <= _T_632_2;
    end
    if (reset) begin
      _T_642_0 <= 1'h0;
    end else begin
      _T_642_0 <= _T_635;
    end
    if (reset) begin
      _T_642_1 <= 1'h0;
    end else begin
      _T_642_1 <= _T_642_0;
    end
    if (reset) begin
      _T_642_2 <= 1'h0;
    end else begin
      _T_642_2 <= _T_642_1;
    end
    if (reset) begin
      _T_642_3 <= 1'h0;
    end else begin
      _T_642_3 <= _T_642_2;
    end
    if (reset) begin
      _T_652_0 <= 1'h0;
    end else begin
      _T_652_0 <= _T_45;
    end
    if (reset) begin
      _T_652_1 <= 1'h0;
    end else begin
      _T_652_1 <= _T_652_0;
    end
    if (reset) begin
      _T_652_2 <= 1'h0;
    end else begin
      _T_652_2 <= _T_652_1;
    end
    if (reset) begin
      _T_652_3 <= 1'h0;
    end else begin
      _T_652_3 <= _T_652_2;
    end
    if (reset) begin
      _T_662_0 <= 1'h0;
    end else begin
      _T_662_0 <= _T_55;
    end
    if (reset) begin
      _T_662_1 <= 1'h0;
    end else begin
      _T_662_1 <= _T_662_0;
    end
    if (reset) begin
      _T_662_2 <= 1'h0;
    end else begin
      _T_662_2 <= _T_662_1;
    end
    if (reset) begin
      _T_662_3 <= 1'h0;
    end else begin
      _T_662_3 <= _T_662_2;
    end
    if (reset) begin
      _T_672_0 <= 1'h0;
    end else begin
      _T_672_0 <= _T_65;
    end
    if (reset) begin
      _T_672_1 <= 1'h0;
    end else begin
      _T_672_1 <= _T_672_0;
    end
    if (reset) begin
      _T_672_2 <= 1'h0;
    end else begin
      _T_672_2 <= _T_672_1;
    end
    if (reset) begin
      _T_672_3 <= 1'h0;
    end else begin
      _T_672_3 <= _T_672_2;
    end
    if (reset) begin
      _T_682_0 <= 1'h0;
    end else begin
      _T_682_0 <= _T_75;
    end
    if (reset) begin
      _T_682_1 <= 1'h0;
    end else begin
      _T_682_1 <= _T_682_0;
    end
    if (reset) begin
      _T_682_2 <= 1'h0;
    end else begin
      _T_682_2 <= _T_682_1;
    end
    if (reset) begin
      _T_682_3 <= 1'h0;
    end else begin
      _T_682_3 <= _T_682_2;
    end
    if (reset) begin
      _T_692_0 <= 1'h0;
    end else begin
      _T_692_0 <= _T_85;
    end
    if (reset) begin
      _T_692_1 <= 1'h0;
    end else begin
      _T_692_1 <= _T_692_0;
    end
    if (reset) begin
      _T_692_2 <= 1'h0;
    end else begin
      _T_692_2 <= _T_692_1;
    end
    if (reset) begin
      _T_692_3 <= 1'h0;
    end else begin
      _T_692_3 <= _T_692_2;
    end
    if (reset) begin
      _T_702_0 <= 1'h0;
    end else begin
      _T_702_0 <= _T_95;
    end
    if (reset) begin
      _T_702_1 <= 1'h0;
    end else begin
      _T_702_1 <= _T_702_0;
    end
    if (reset) begin
      _T_702_2 <= 1'h0;
    end else begin
      _T_702_2 <= _T_702_1;
    end
    if (reset) begin
      _T_702_3 <= 1'h0;
    end else begin
      _T_702_3 <= _T_702_2;
    end
    if (reset) begin
      _T_712_0 <= 1'h0;
    end else begin
      _T_712_0 <= _T_105;
    end
    if (reset) begin
      _T_712_1 <= 1'h0;
    end else begin
      _T_712_1 <= _T_712_0;
    end
    if (reset) begin
      _T_712_2 <= 1'h0;
    end else begin
      _T_712_2 <= _T_712_1;
    end
    if (reset) begin
      _T_712_3 <= 1'h0;
    end else begin
      _T_712_3 <= _T_712_2;
    end
    if (reset) begin
      _T_722_0 <= 1'h0;
    end else begin
      _T_722_0 <= _T_115;
    end
    if (reset) begin
      _T_722_1 <= 1'h0;
    end else begin
      _T_722_1 <= _T_722_0;
    end
    if (reset) begin
      _T_722_2 <= 1'h0;
    end else begin
      _T_722_2 <= _T_722_1;
    end
    if (reset) begin
      _T_722_3 <= 1'h0;
    end else begin
      _T_722_3 <= _T_722_2;
    end
    if (reset) begin
      _T_732_0 <= 1'h0;
    end else begin
      _T_732_0 <= _T_125;
    end
    if (reset) begin
      _T_732_1 <= 1'h0;
    end else begin
      _T_732_1 <= _T_732_0;
    end
    if (reset) begin
      _T_732_2 <= 1'h0;
    end else begin
      _T_732_2 <= _T_732_1;
    end
    if (reset) begin
      _T_732_3 <= 1'h0;
    end else begin
      _T_732_3 <= _T_732_2;
    end
    if (reset) begin
      _T_742_0 <= 1'h0;
    end else begin
      _T_742_0 <= _T_135;
    end
    if (reset) begin
      _T_742_1 <= 1'h0;
    end else begin
      _T_742_1 <= _T_742_0;
    end
    if (reset) begin
      _T_742_2 <= 1'h0;
    end else begin
      _T_742_2 <= _T_742_1;
    end
    if (reset) begin
      _T_742_3 <= 1'h0;
    end else begin
      _T_742_3 <= _T_742_2;
    end
    if (reset) begin
      _T_752_0 <= 1'h0;
    end else begin
      _T_752_0 <= _T_145;
    end
    if (reset) begin
      _T_752_1 <= 1'h0;
    end else begin
      _T_752_1 <= _T_752_0;
    end
    if (reset) begin
      _T_752_2 <= 1'h0;
    end else begin
      _T_752_2 <= _T_752_1;
    end
    if (reset) begin
      _T_752_3 <= 1'h0;
    end else begin
      _T_752_3 <= _T_752_2;
    end
    if (reset) begin
      _T_762_0 <= 1'h0;
    end else begin
      _T_762_0 <= _T_155;
    end
    if (reset) begin
      _T_762_1 <= 1'h0;
    end else begin
      _T_762_1 <= _T_762_0;
    end
    if (reset) begin
      _T_762_2 <= 1'h0;
    end else begin
      _T_762_2 <= _T_762_1;
    end
    if (reset) begin
      _T_762_3 <= 1'h0;
    end else begin
      _T_762_3 <= _T_762_2;
    end
    if (reset) begin
      _T_772_0 <= 1'h0;
    end else begin
      _T_772_0 <= _T_315;
    end
    if (reset) begin
      _T_772_1 <= 1'h0;
    end else begin
      _T_772_1 <= _T_772_0;
    end
    if (reset) begin
      _T_772_2 <= 1'h0;
    end else begin
      _T_772_2 <= _T_772_1;
    end
    if (reset) begin
      _T_772_3 <= 1'h0;
    end else begin
      _T_772_3 <= _T_772_2;
    end
    if (reset) begin
      _T_782_0 <= 1'h0;
    end else begin
      _T_782_0 <= _T_475;
    end
    if (reset) begin
      _T_782_1 <= 1'h0;
    end else begin
      _T_782_1 <= _T_782_0;
    end
    if (reset) begin
      _T_782_2 <= 1'h0;
    end else begin
      _T_782_2 <= _T_782_1;
    end
    if (reset) begin
      _T_782_3 <= 1'h0;
    end else begin
      _T_782_3 <= _T_782_2;
    end
    if (reset) begin
      _T_792_0 <= 1'h0;
    end else begin
      _T_792_0 <= _T_635;
    end
    if (reset) begin
      _T_792_1 <= 1'h0;
    end else begin
      _T_792_1 <= _T_792_0;
    end
    if (reset) begin
      _T_792_2 <= 1'h0;
    end else begin
      _T_792_2 <= _T_792_1;
    end
    if (reset) begin
      _T_792_3 <= 1'h0;
    end else begin
      _T_792_3 <= _T_792_2;
    end
    if (reset) begin
      _T_802_0 <= 1'h0;
    end else begin
      _T_802_0 <= _T_795;
    end
    if (reset) begin
      _T_802_1 <= 1'h0;
    end else begin
      _T_802_1 <= _T_802_0;
    end
    if (reset) begin
      _T_802_2 <= 1'h0;
    end else begin
      _T_802_2 <= _T_802_1;
    end
    if (reset) begin
      _T_802_3 <= 1'h0;
    end else begin
      _T_802_3 <= _T_802_2;
    end
    if (reset) begin
      _T_812_0 <= 1'h0;
    end else begin
      _T_812_0 <= _T_55;
    end
    if (reset) begin
      _T_812_1 <= 1'h0;
    end else begin
      _T_812_1 <= _T_812_0;
    end
    if (reset) begin
      _T_812_2 <= 1'h0;
    end else begin
      _T_812_2 <= _T_812_1;
    end
    if (reset) begin
      _T_812_3 <= 1'h0;
    end else begin
      _T_812_3 <= _T_812_2;
    end
    if (reset) begin
      _T_822_0 <= 1'h0;
    end else begin
      _T_822_0 <= _T_65;
    end
    if (reset) begin
      _T_822_1 <= 1'h0;
    end else begin
      _T_822_1 <= _T_822_0;
    end
    if (reset) begin
      _T_822_2 <= 1'h0;
    end else begin
      _T_822_2 <= _T_822_1;
    end
    if (reset) begin
      _T_822_3 <= 1'h0;
    end else begin
      _T_822_3 <= _T_822_2;
    end
    if (reset) begin
      _T_832_0 <= 1'h0;
    end else begin
      _T_832_0 <= _T_75;
    end
    if (reset) begin
      _T_832_1 <= 1'h0;
    end else begin
      _T_832_1 <= _T_832_0;
    end
    if (reset) begin
      _T_832_2 <= 1'h0;
    end else begin
      _T_832_2 <= _T_832_1;
    end
    if (reset) begin
      _T_832_3 <= 1'h0;
    end else begin
      _T_832_3 <= _T_832_2;
    end
    if (reset) begin
      _T_842_0 <= 1'h0;
    end else begin
      _T_842_0 <= _T_85;
    end
    if (reset) begin
      _T_842_1 <= 1'h0;
    end else begin
      _T_842_1 <= _T_842_0;
    end
    if (reset) begin
      _T_842_2 <= 1'h0;
    end else begin
      _T_842_2 <= _T_842_1;
    end
    if (reset) begin
      _T_842_3 <= 1'h0;
    end else begin
      _T_842_3 <= _T_842_2;
    end
    if (reset) begin
      _T_852_0 <= 1'h0;
    end else begin
      _T_852_0 <= _T_95;
    end
    if (reset) begin
      _T_852_1 <= 1'h0;
    end else begin
      _T_852_1 <= _T_852_0;
    end
    if (reset) begin
      _T_852_2 <= 1'h0;
    end else begin
      _T_852_2 <= _T_852_1;
    end
    if (reset) begin
      _T_852_3 <= 1'h0;
    end else begin
      _T_852_3 <= _T_852_2;
    end
    if (reset) begin
      _T_862_0 <= 1'h0;
    end else begin
      _T_862_0 <= _T_105;
    end
    if (reset) begin
      _T_862_1 <= 1'h0;
    end else begin
      _T_862_1 <= _T_862_0;
    end
    if (reset) begin
      _T_862_2 <= 1'h0;
    end else begin
      _T_862_2 <= _T_862_1;
    end
    if (reset) begin
      _T_862_3 <= 1'h0;
    end else begin
      _T_862_3 <= _T_862_2;
    end
    if (reset) begin
      _T_872_0 <= 1'h0;
    end else begin
      _T_872_0 <= _T_115;
    end
    if (reset) begin
      _T_872_1 <= 1'h0;
    end else begin
      _T_872_1 <= _T_872_0;
    end
    if (reset) begin
      _T_872_2 <= 1'h0;
    end else begin
      _T_872_2 <= _T_872_1;
    end
    if (reset) begin
      _T_872_3 <= 1'h0;
    end else begin
      _T_872_3 <= _T_872_2;
    end
    if (reset) begin
      _T_882_0 <= 1'h0;
    end else begin
      _T_882_0 <= _T_125;
    end
    if (reset) begin
      _T_882_1 <= 1'h0;
    end else begin
      _T_882_1 <= _T_882_0;
    end
    if (reset) begin
      _T_882_2 <= 1'h0;
    end else begin
      _T_882_2 <= _T_882_1;
    end
    if (reset) begin
      _T_882_3 <= 1'h0;
    end else begin
      _T_882_3 <= _T_882_2;
    end
    if (reset) begin
      _T_892_0 <= 1'h0;
    end else begin
      _T_892_0 <= _T_135;
    end
    if (reset) begin
      _T_892_1 <= 1'h0;
    end else begin
      _T_892_1 <= _T_892_0;
    end
    if (reset) begin
      _T_892_2 <= 1'h0;
    end else begin
      _T_892_2 <= _T_892_1;
    end
    if (reset) begin
      _T_892_3 <= 1'h0;
    end else begin
      _T_892_3 <= _T_892_2;
    end
    if (reset) begin
      _T_902_0 <= 1'h0;
    end else begin
      _T_902_0 <= _T_145;
    end
    if (reset) begin
      _T_902_1 <= 1'h0;
    end else begin
      _T_902_1 <= _T_902_0;
    end
    if (reset) begin
      _T_902_2 <= 1'h0;
    end else begin
      _T_902_2 <= _T_902_1;
    end
    if (reset) begin
      _T_902_3 <= 1'h0;
    end else begin
      _T_902_3 <= _T_902_2;
    end
    if (reset) begin
      _T_912_0 <= 1'h0;
    end else begin
      _T_912_0 <= _T_155;
    end
    if (reset) begin
      _T_912_1 <= 1'h0;
    end else begin
      _T_912_1 <= _T_912_0;
    end
    if (reset) begin
      _T_912_2 <= 1'h0;
    end else begin
      _T_912_2 <= _T_912_1;
    end
    if (reset) begin
      _T_912_3 <= 1'h0;
    end else begin
      _T_912_3 <= _T_912_2;
    end
    if (reset) begin
      _T_922_0 <= 1'h0;
    end else begin
      _T_922_0 <= _T_315;
    end
    if (reset) begin
      _T_922_1 <= 1'h0;
    end else begin
      _T_922_1 <= _T_922_0;
    end
    if (reset) begin
      _T_922_2 <= 1'h0;
    end else begin
      _T_922_2 <= _T_922_1;
    end
    if (reset) begin
      _T_922_3 <= 1'h0;
    end else begin
      _T_922_3 <= _T_922_2;
    end
    if (reset) begin
      _T_932_0 <= 1'h0;
    end else begin
      _T_932_0 <= _T_475;
    end
    if (reset) begin
      _T_932_1 <= 1'h0;
    end else begin
      _T_932_1 <= _T_932_0;
    end
    if (reset) begin
      _T_932_2 <= 1'h0;
    end else begin
      _T_932_2 <= _T_932_1;
    end
    if (reset) begin
      _T_932_3 <= 1'h0;
    end else begin
      _T_932_3 <= _T_932_2;
    end
    if (reset) begin
      _T_942_0 <= 1'h0;
    end else begin
      _T_942_0 <= _T_635;
    end
    if (reset) begin
      _T_942_1 <= 1'h0;
    end else begin
      _T_942_1 <= _T_942_0;
    end
    if (reset) begin
      _T_942_2 <= 1'h0;
    end else begin
      _T_942_2 <= _T_942_1;
    end
    if (reset) begin
      _T_942_3 <= 1'h0;
    end else begin
      _T_942_3 <= _T_942_2;
    end
    if (reset) begin
      _T_952_0 <= 1'h0;
    end else begin
      _T_952_0 <= _T_795;
    end
    if (reset) begin
      _T_952_1 <= 1'h0;
    end else begin
      _T_952_1 <= _T_952_0;
    end
    if (reset) begin
      _T_952_2 <= 1'h0;
    end else begin
      _T_952_2 <= _T_952_1;
    end
    if (reset) begin
      _T_952_3 <= 1'h0;
    end else begin
      _T_952_3 <= _T_952_2;
    end
    if (reset) begin
      _T_962_0 <= 1'h0;
    end else begin
      _T_962_0 <= _T_955;
    end
    if (reset) begin
      _T_962_1 <= 1'h0;
    end else begin
      _T_962_1 <= _T_962_0;
    end
    if (reset) begin
      _T_962_2 <= 1'h0;
    end else begin
      _T_962_2 <= _T_962_1;
    end
    if (reset) begin
      _T_962_3 <= 1'h0;
    end else begin
      _T_962_3 <= _T_962_2;
    end
    if (reset) begin
      _T_972_0 <= 1'h0;
    end else begin
      _T_972_0 <= _T_65;
    end
    if (reset) begin
      _T_972_1 <= 1'h0;
    end else begin
      _T_972_1 <= _T_972_0;
    end
    if (reset) begin
      _T_972_2 <= 1'h0;
    end else begin
      _T_972_2 <= _T_972_1;
    end
    if (reset) begin
      _T_972_3 <= 1'h0;
    end else begin
      _T_972_3 <= _T_972_2;
    end
    if (reset) begin
      _T_982_0 <= 1'h0;
    end else begin
      _T_982_0 <= _T_75;
    end
    if (reset) begin
      _T_982_1 <= 1'h0;
    end else begin
      _T_982_1 <= _T_982_0;
    end
    if (reset) begin
      _T_982_2 <= 1'h0;
    end else begin
      _T_982_2 <= _T_982_1;
    end
    if (reset) begin
      _T_982_3 <= 1'h0;
    end else begin
      _T_982_3 <= _T_982_2;
    end
    if (reset) begin
      _T_992_0 <= 1'h0;
    end else begin
      _T_992_0 <= _T_85;
    end
    if (reset) begin
      _T_992_1 <= 1'h0;
    end else begin
      _T_992_1 <= _T_992_0;
    end
    if (reset) begin
      _T_992_2 <= 1'h0;
    end else begin
      _T_992_2 <= _T_992_1;
    end
    if (reset) begin
      _T_992_3 <= 1'h0;
    end else begin
      _T_992_3 <= _T_992_2;
    end
    if (reset) begin
      _T_1002_0 <= 1'h0;
    end else begin
      _T_1002_0 <= _T_95;
    end
    if (reset) begin
      _T_1002_1 <= 1'h0;
    end else begin
      _T_1002_1 <= _T_1002_0;
    end
    if (reset) begin
      _T_1002_2 <= 1'h0;
    end else begin
      _T_1002_2 <= _T_1002_1;
    end
    if (reset) begin
      _T_1002_3 <= 1'h0;
    end else begin
      _T_1002_3 <= _T_1002_2;
    end
    if (reset) begin
      _T_1012_0 <= 1'h0;
    end else begin
      _T_1012_0 <= _T_105;
    end
    if (reset) begin
      _T_1012_1 <= 1'h0;
    end else begin
      _T_1012_1 <= _T_1012_0;
    end
    if (reset) begin
      _T_1012_2 <= 1'h0;
    end else begin
      _T_1012_2 <= _T_1012_1;
    end
    if (reset) begin
      _T_1012_3 <= 1'h0;
    end else begin
      _T_1012_3 <= _T_1012_2;
    end
    if (reset) begin
      _T_1022_0 <= 1'h0;
    end else begin
      _T_1022_0 <= _T_115;
    end
    if (reset) begin
      _T_1022_1 <= 1'h0;
    end else begin
      _T_1022_1 <= _T_1022_0;
    end
    if (reset) begin
      _T_1022_2 <= 1'h0;
    end else begin
      _T_1022_2 <= _T_1022_1;
    end
    if (reset) begin
      _T_1022_3 <= 1'h0;
    end else begin
      _T_1022_3 <= _T_1022_2;
    end
    if (reset) begin
      _T_1032_0 <= 1'h0;
    end else begin
      _T_1032_0 <= _T_125;
    end
    if (reset) begin
      _T_1032_1 <= 1'h0;
    end else begin
      _T_1032_1 <= _T_1032_0;
    end
    if (reset) begin
      _T_1032_2 <= 1'h0;
    end else begin
      _T_1032_2 <= _T_1032_1;
    end
    if (reset) begin
      _T_1032_3 <= 1'h0;
    end else begin
      _T_1032_3 <= _T_1032_2;
    end
    if (reset) begin
      _T_1042_0 <= 1'h0;
    end else begin
      _T_1042_0 <= _T_135;
    end
    if (reset) begin
      _T_1042_1 <= 1'h0;
    end else begin
      _T_1042_1 <= _T_1042_0;
    end
    if (reset) begin
      _T_1042_2 <= 1'h0;
    end else begin
      _T_1042_2 <= _T_1042_1;
    end
    if (reset) begin
      _T_1042_3 <= 1'h0;
    end else begin
      _T_1042_3 <= _T_1042_2;
    end
    if (reset) begin
      _T_1052_0 <= 1'h0;
    end else begin
      _T_1052_0 <= _T_145;
    end
    if (reset) begin
      _T_1052_1 <= 1'h0;
    end else begin
      _T_1052_1 <= _T_1052_0;
    end
    if (reset) begin
      _T_1052_2 <= 1'h0;
    end else begin
      _T_1052_2 <= _T_1052_1;
    end
    if (reset) begin
      _T_1052_3 <= 1'h0;
    end else begin
      _T_1052_3 <= _T_1052_2;
    end
    if (reset) begin
      _T_1062_0 <= 1'h0;
    end else begin
      _T_1062_0 <= _T_155;
    end
    if (reset) begin
      _T_1062_1 <= 1'h0;
    end else begin
      _T_1062_1 <= _T_1062_0;
    end
    if (reset) begin
      _T_1062_2 <= 1'h0;
    end else begin
      _T_1062_2 <= _T_1062_1;
    end
    if (reset) begin
      _T_1062_3 <= 1'h0;
    end else begin
      _T_1062_3 <= _T_1062_2;
    end
    if (reset) begin
      _T_1072_0 <= 1'h0;
    end else begin
      _T_1072_0 <= _T_315;
    end
    if (reset) begin
      _T_1072_1 <= 1'h0;
    end else begin
      _T_1072_1 <= _T_1072_0;
    end
    if (reset) begin
      _T_1072_2 <= 1'h0;
    end else begin
      _T_1072_2 <= _T_1072_1;
    end
    if (reset) begin
      _T_1072_3 <= 1'h0;
    end else begin
      _T_1072_3 <= _T_1072_2;
    end
    if (reset) begin
      _T_1082_0 <= 1'h0;
    end else begin
      _T_1082_0 <= _T_475;
    end
    if (reset) begin
      _T_1082_1 <= 1'h0;
    end else begin
      _T_1082_1 <= _T_1082_0;
    end
    if (reset) begin
      _T_1082_2 <= 1'h0;
    end else begin
      _T_1082_2 <= _T_1082_1;
    end
    if (reset) begin
      _T_1082_3 <= 1'h0;
    end else begin
      _T_1082_3 <= _T_1082_2;
    end
    if (reset) begin
      _T_1092_0 <= 1'h0;
    end else begin
      _T_1092_0 <= _T_635;
    end
    if (reset) begin
      _T_1092_1 <= 1'h0;
    end else begin
      _T_1092_1 <= _T_1092_0;
    end
    if (reset) begin
      _T_1092_2 <= 1'h0;
    end else begin
      _T_1092_2 <= _T_1092_1;
    end
    if (reset) begin
      _T_1092_3 <= 1'h0;
    end else begin
      _T_1092_3 <= _T_1092_2;
    end
    if (reset) begin
      _T_1102_0 <= 1'h0;
    end else begin
      _T_1102_0 <= _T_795;
    end
    if (reset) begin
      _T_1102_1 <= 1'h0;
    end else begin
      _T_1102_1 <= _T_1102_0;
    end
    if (reset) begin
      _T_1102_2 <= 1'h0;
    end else begin
      _T_1102_2 <= _T_1102_1;
    end
    if (reset) begin
      _T_1102_3 <= 1'h0;
    end else begin
      _T_1102_3 <= _T_1102_2;
    end
    if (reset) begin
      _T_1112_0 <= 1'h0;
    end else begin
      _T_1112_0 <= _T_955;
    end
    if (reset) begin
      _T_1112_1 <= 1'h0;
    end else begin
      _T_1112_1 <= _T_1112_0;
    end
    if (reset) begin
      _T_1112_2 <= 1'h0;
    end else begin
      _T_1112_2 <= _T_1112_1;
    end
    if (reset) begin
      _T_1112_3 <= 1'h0;
    end else begin
      _T_1112_3 <= _T_1112_2;
    end
    if (reset) begin
      _T_1122_0 <= 1'h0;
    end else begin
      _T_1122_0 <= _T_1115;
    end
    if (reset) begin
      _T_1122_1 <= 1'h0;
    end else begin
      _T_1122_1 <= _T_1122_0;
    end
    if (reset) begin
      _T_1122_2 <= 1'h0;
    end else begin
      _T_1122_2 <= _T_1122_1;
    end
    if (reset) begin
      _T_1122_3 <= 1'h0;
    end else begin
      _T_1122_3 <= _T_1122_2;
    end
    if (reset) begin
      _T_1132_0 <= 1'h0;
    end else begin
      _T_1132_0 <= _T_75;
    end
    if (reset) begin
      _T_1132_1 <= 1'h0;
    end else begin
      _T_1132_1 <= _T_1132_0;
    end
    if (reset) begin
      _T_1132_2 <= 1'h0;
    end else begin
      _T_1132_2 <= _T_1132_1;
    end
    if (reset) begin
      _T_1132_3 <= 1'h0;
    end else begin
      _T_1132_3 <= _T_1132_2;
    end
    if (reset) begin
      _T_1142_0 <= 1'h0;
    end else begin
      _T_1142_0 <= _T_85;
    end
    if (reset) begin
      _T_1142_1 <= 1'h0;
    end else begin
      _T_1142_1 <= _T_1142_0;
    end
    if (reset) begin
      _T_1142_2 <= 1'h0;
    end else begin
      _T_1142_2 <= _T_1142_1;
    end
    if (reset) begin
      _T_1142_3 <= 1'h0;
    end else begin
      _T_1142_3 <= _T_1142_2;
    end
    if (reset) begin
      _T_1152_0 <= 1'h0;
    end else begin
      _T_1152_0 <= _T_95;
    end
    if (reset) begin
      _T_1152_1 <= 1'h0;
    end else begin
      _T_1152_1 <= _T_1152_0;
    end
    if (reset) begin
      _T_1152_2 <= 1'h0;
    end else begin
      _T_1152_2 <= _T_1152_1;
    end
    if (reset) begin
      _T_1152_3 <= 1'h0;
    end else begin
      _T_1152_3 <= _T_1152_2;
    end
    if (reset) begin
      _T_1162_0 <= 1'h0;
    end else begin
      _T_1162_0 <= _T_105;
    end
    if (reset) begin
      _T_1162_1 <= 1'h0;
    end else begin
      _T_1162_1 <= _T_1162_0;
    end
    if (reset) begin
      _T_1162_2 <= 1'h0;
    end else begin
      _T_1162_2 <= _T_1162_1;
    end
    if (reset) begin
      _T_1162_3 <= 1'h0;
    end else begin
      _T_1162_3 <= _T_1162_2;
    end
    if (reset) begin
      _T_1172_0 <= 1'h0;
    end else begin
      _T_1172_0 <= _T_115;
    end
    if (reset) begin
      _T_1172_1 <= 1'h0;
    end else begin
      _T_1172_1 <= _T_1172_0;
    end
    if (reset) begin
      _T_1172_2 <= 1'h0;
    end else begin
      _T_1172_2 <= _T_1172_1;
    end
    if (reset) begin
      _T_1172_3 <= 1'h0;
    end else begin
      _T_1172_3 <= _T_1172_2;
    end
    if (reset) begin
      _T_1182_0 <= 1'h0;
    end else begin
      _T_1182_0 <= _T_125;
    end
    if (reset) begin
      _T_1182_1 <= 1'h0;
    end else begin
      _T_1182_1 <= _T_1182_0;
    end
    if (reset) begin
      _T_1182_2 <= 1'h0;
    end else begin
      _T_1182_2 <= _T_1182_1;
    end
    if (reset) begin
      _T_1182_3 <= 1'h0;
    end else begin
      _T_1182_3 <= _T_1182_2;
    end
    if (reset) begin
      _T_1192_0 <= 1'h0;
    end else begin
      _T_1192_0 <= _T_135;
    end
    if (reset) begin
      _T_1192_1 <= 1'h0;
    end else begin
      _T_1192_1 <= _T_1192_0;
    end
    if (reset) begin
      _T_1192_2 <= 1'h0;
    end else begin
      _T_1192_2 <= _T_1192_1;
    end
    if (reset) begin
      _T_1192_3 <= 1'h0;
    end else begin
      _T_1192_3 <= _T_1192_2;
    end
    if (reset) begin
      _T_1202_0 <= 1'h0;
    end else begin
      _T_1202_0 <= _T_145;
    end
    if (reset) begin
      _T_1202_1 <= 1'h0;
    end else begin
      _T_1202_1 <= _T_1202_0;
    end
    if (reset) begin
      _T_1202_2 <= 1'h0;
    end else begin
      _T_1202_2 <= _T_1202_1;
    end
    if (reset) begin
      _T_1202_3 <= 1'h0;
    end else begin
      _T_1202_3 <= _T_1202_2;
    end
    if (reset) begin
      _T_1212_0 <= 1'h0;
    end else begin
      _T_1212_0 <= _T_155;
    end
    if (reset) begin
      _T_1212_1 <= 1'h0;
    end else begin
      _T_1212_1 <= _T_1212_0;
    end
    if (reset) begin
      _T_1212_2 <= 1'h0;
    end else begin
      _T_1212_2 <= _T_1212_1;
    end
    if (reset) begin
      _T_1212_3 <= 1'h0;
    end else begin
      _T_1212_3 <= _T_1212_2;
    end
    if (reset) begin
      _T_1222_0 <= 1'h0;
    end else begin
      _T_1222_0 <= _T_315;
    end
    if (reset) begin
      _T_1222_1 <= 1'h0;
    end else begin
      _T_1222_1 <= _T_1222_0;
    end
    if (reset) begin
      _T_1222_2 <= 1'h0;
    end else begin
      _T_1222_2 <= _T_1222_1;
    end
    if (reset) begin
      _T_1222_3 <= 1'h0;
    end else begin
      _T_1222_3 <= _T_1222_2;
    end
    if (reset) begin
      _T_1232_0 <= 1'h0;
    end else begin
      _T_1232_0 <= _T_475;
    end
    if (reset) begin
      _T_1232_1 <= 1'h0;
    end else begin
      _T_1232_1 <= _T_1232_0;
    end
    if (reset) begin
      _T_1232_2 <= 1'h0;
    end else begin
      _T_1232_2 <= _T_1232_1;
    end
    if (reset) begin
      _T_1232_3 <= 1'h0;
    end else begin
      _T_1232_3 <= _T_1232_2;
    end
    if (reset) begin
      _T_1242_0 <= 1'h0;
    end else begin
      _T_1242_0 <= _T_635;
    end
    if (reset) begin
      _T_1242_1 <= 1'h0;
    end else begin
      _T_1242_1 <= _T_1242_0;
    end
    if (reset) begin
      _T_1242_2 <= 1'h0;
    end else begin
      _T_1242_2 <= _T_1242_1;
    end
    if (reset) begin
      _T_1242_3 <= 1'h0;
    end else begin
      _T_1242_3 <= _T_1242_2;
    end
    if (reset) begin
      _T_1252_0 <= 1'h0;
    end else begin
      _T_1252_0 <= _T_795;
    end
    if (reset) begin
      _T_1252_1 <= 1'h0;
    end else begin
      _T_1252_1 <= _T_1252_0;
    end
    if (reset) begin
      _T_1252_2 <= 1'h0;
    end else begin
      _T_1252_2 <= _T_1252_1;
    end
    if (reset) begin
      _T_1252_3 <= 1'h0;
    end else begin
      _T_1252_3 <= _T_1252_2;
    end
    if (reset) begin
      _T_1262_0 <= 1'h0;
    end else begin
      _T_1262_0 <= _T_955;
    end
    if (reset) begin
      _T_1262_1 <= 1'h0;
    end else begin
      _T_1262_1 <= _T_1262_0;
    end
    if (reset) begin
      _T_1262_2 <= 1'h0;
    end else begin
      _T_1262_2 <= _T_1262_1;
    end
    if (reset) begin
      _T_1262_3 <= 1'h0;
    end else begin
      _T_1262_3 <= _T_1262_2;
    end
    if (reset) begin
      _T_1272_0 <= 1'h0;
    end else begin
      _T_1272_0 <= _T_1115;
    end
    if (reset) begin
      _T_1272_1 <= 1'h0;
    end else begin
      _T_1272_1 <= _T_1272_0;
    end
    if (reset) begin
      _T_1272_2 <= 1'h0;
    end else begin
      _T_1272_2 <= _T_1272_1;
    end
    if (reset) begin
      _T_1272_3 <= 1'h0;
    end else begin
      _T_1272_3 <= _T_1272_2;
    end
    if (reset) begin
      _T_1282_0 <= 1'h0;
    end else begin
      _T_1282_0 <= _T_1275;
    end
    if (reset) begin
      _T_1282_1 <= 1'h0;
    end else begin
      _T_1282_1 <= _T_1282_0;
    end
    if (reset) begin
      _T_1282_2 <= 1'h0;
    end else begin
      _T_1282_2 <= _T_1282_1;
    end
    if (reset) begin
      _T_1282_3 <= 1'h0;
    end else begin
      _T_1282_3 <= _T_1282_2;
    end
    if (reset) begin
      _T_1292_0 <= 1'h0;
    end else begin
      _T_1292_0 <= _T_85;
    end
    if (reset) begin
      _T_1292_1 <= 1'h0;
    end else begin
      _T_1292_1 <= _T_1292_0;
    end
    if (reset) begin
      _T_1292_2 <= 1'h0;
    end else begin
      _T_1292_2 <= _T_1292_1;
    end
    if (reset) begin
      _T_1292_3 <= 1'h0;
    end else begin
      _T_1292_3 <= _T_1292_2;
    end
    if (reset) begin
      _T_1302_0 <= 1'h0;
    end else begin
      _T_1302_0 <= _T_95;
    end
    if (reset) begin
      _T_1302_1 <= 1'h0;
    end else begin
      _T_1302_1 <= _T_1302_0;
    end
    if (reset) begin
      _T_1302_2 <= 1'h0;
    end else begin
      _T_1302_2 <= _T_1302_1;
    end
    if (reset) begin
      _T_1302_3 <= 1'h0;
    end else begin
      _T_1302_3 <= _T_1302_2;
    end
    if (reset) begin
      _T_1312_0 <= 1'h0;
    end else begin
      _T_1312_0 <= _T_105;
    end
    if (reset) begin
      _T_1312_1 <= 1'h0;
    end else begin
      _T_1312_1 <= _T_1312_0;
    end
    if (reset) begin
      _T_1312_2 <= 1'h0;
    end else begin
      _T_1312_2 <= _T_1312_1;
    end
    if (reset) begin
      _T_1312_3 <= 1'h0;
    end else begin
      _T_1312_3 <= _T_1312_2;
    end
    if (reset) begin
      _T_1322_0 <= 1'h0;
    end else begin
      _T_1322_0 <= _T_115;
    end
    if (reset) begin
      _T_1322_1 <= 1'h0;
    end else begin
      _T_1322_1 <= _T_1322_0;
    end
    if (reset) begin
      _T_1322_2 <= 1'h0;
    end else begin
      _T_1322_2 <= _T_1322_1;
    end
    if (reset) begin
      _T_1322_3 <= 1'h0;
    end else begin
      _T_1322_3 <= _T_1322_2;
    end
    if (reset) begin
      _T_1332_0 <= 1'h0;
    end else begin
      _T_1332_0 <= _T_125;
    end
    if (reset) begin
      _T_1332_1 <= 1'h0;
    end else begin
      _T_1332_1 <= _T_1332_0;
    end
    if (reset) begin
      _T_1332_2 <= 1'h0;
    end else begin
      _T_1332_2 <= _T_1332_1;
    end
    if (reset) begin
      _T_1332_3 <= 1'h0;
    end else begin
      _T_1332_3 <= _T_1332_2;
    end
    if (reset) begin
      _T_1342_0 <= 1'h0;
    end else begin
      _T_1342_0 <= _T_135;
    end
    if (reset) begin
      _T_1342_1 <= 1'h0;
    end else begin
      _T_1342_1 <= _T_1342_0;
    end
    if (reset) begin
      _T_1342_2 <= 1'h0;
    end else begin
      _T_1342_2 <= _T_1342_1;
    end
    if (reset) begin
      _T_1342_3 <= 1'h0;
    end else begin
      _T_1342_3 <= _T_1342_2;
    end
    if (reset) begin
      _T_1352_0 <= 1'h0;
    end else begin
      _T_1352_0 <= _T_145;
    end
    if (reset) begin
      _T_1352_1 <= 1'h0;
    end else begin
      _T_1352_1 <= _T_1352_0;
    end
    if (reset) begin
      _T_1352_2 <= 1'h0;
    end else begin
      _T_1352_2 <= _T_1352_1;
    end
    if (reset) begin
      _T_1352_3 <= 1'h0;
    end else begin
      _T_1352_3 <= _T_1352_2;
    end
    if (reset) begin
      _T_1362_0 <= 1'h0;
    end else begin
      _T_1362_0 <= _T_155;
    end
    if (reset) begin
      _T_1362_1 <= 1'h0;
    end else begin
      _T_1362_1 <= _T_1362_0;
    end
    if (reset) begin
      _T_1362_2 <= 1'h0;
    end else begin
      _T_1362_2 <= _T_1362_1;
    end
    if (reset) begin
      _T_1362_3 <= 1'h0;
    end else begin
      _T_1362_3 <= _T_1362_2;
    end
    if (reset) begin
      _T_1372_0 <= 1'h0;
    end else begin
      _T_1372_0 <= _T_315;
    end
    if (reset) begin
      _T_1372_1 <= 1'h0;
    end else begin
      _T_1372_1 <= _T_1372_0;
    end
    if (reset) begin
      _T_1372_2 <= 1'h0;
    end else begin
      _T_1372_2 <= _T_1372_1;
    end
    if (reset) begin
      _T_1372_3 <= 1'h0;
    end else begin
      _T_1372_3 <= _T_1372_2;
    end
    if (reset) begin
      _T_1382_0 <= 1'h0;
    end else begin
      _T_1382_0 <= _T_475;
    end
    if (reset) begin
      _T_1382_1 <= 1'h0;
    end else begin
      _T_1382_1 <= _T_1382_0;
    end
    if (reset) begin
      _T_1382_2 <= 1'h0;
    end else begin
      _T_1382_2 <= _T_1382_1;
    end
    if (reset) begin
      _T_1382_3 <= 1'h0;
    end else begin
      _T_1382_3 <= _T_1382_2;
    end
    if (reset) begin
      _T_1392_0 <= 1'h0;
    end else begin
      _T_1392_0 <= _T_635;
    end
    if (reset) begin
      _T_1392_1 <= 1'h0;
    end else begin
      _T_1392_1 <= _T_1392_0;
    end
    if (reset) begin
      _T_1392_2 <= 1'h0;
    end else begin
      _T_1392_2 <= _T_1392_1;
    end
    if (reset) begin
      _T_1392_3 <= 1'h0;
    end else begin
      _T_1392_3 <= _T_1392_2;
    end
    if (reset) begin
      _T_1402_0 <= 1'h0;
    end else begin
      _T_1402_0 <= _T_795;
    end
    if (reset) begin
      _T_1402_1 <= 1'h0;
    end else begin
      _T_1402_1 <= _T_1402_0;
    end
    if (reset) begin
      _T_1402_2 <= 1'h0;
    end else begin
      _T_1402_2 <= _T_1402_1;
    end
    if (reset) begin
      _T_1402_3 <= 1'h0;
    end else begin
      _T_1402_3 <= _T_1402_2;
    end
    if (reset) begin
      _T_1412_0 <= 1'h0;
    end else begin
      _T_1412_0 <= _T_955;
    end
    if (reset) begin
      _T_1412_1 <= 1'h0;
    end else begin
      _T_1412_1 <= _T_1412_0;
    end
    if (reset) begin
      _T_1412_2 <= 1'h0;
    end else begin
      _T_1412_2 <= _T_1412_1;
    end
    if (reset) begin
      _T_1412_3 <= 1'h0;
    end else begin
      _T_1412_3 <= _T_1412_2;
    end
    if (reset) begin
      _T_1422_0 <= 1'h0;
    end else begin
      _T_1422_0 <= _T_1115;
    end
    if (reset) begin
      _T_1422_1 <= 1'h0;
    end else begin
      _T_1422_1 <= _T_1422_0;
    end
    if (reset) begin
      _T_1422_2 <= 1'h0;
    end else begin
      _T_1422_2 <= _T_1422_1;
    end
    if (reset) begin
      _T_1422_3 <= 1'h0;
    end else begin
      _T_1422_3 <= _T_1422_2;
    end
    if (reset) begin
      _T_1432_0 <= 1'h0;
    end else begin
      _T_1432_0 <= _T_1275;
    end
    if (reset) begin
      _T_1432_1 <= 1'h0;
    end else begin
      _T_1432_1 <= _T_1432_0;
    end
    if (reset) begin
      _T_1432_2 <= 1'h0;
    end else begin
      _T_1432_2 <= _T_1432_1;
    end
    if (reset) begin
      _T_1432_3 <= 1'h0;
    end else begin
      _T_1432_3 <= _T_1432_2;
    end
    if (reset) begin
      _T_1442_0 <= 1'h0;
    end else begin
      _T_1442_0 <= _T_1435;
    end
    if (reset) begin
      _T_1442_1 <= 1'h0;
    end else begin
      _T_1442_1 <= _T_1442_0;
    end
    if (reset) begin
      _T_1442_2 <= 1'h0;
    end else begin
      _T_1442_2 <= _T_1442_1;
    end
    if (reset) begin
      _T_1442_3 <= 1'h0;
    end else begin
      _T_1442_3 <= _T_1442_2;
    end
    if (reset) begin
      _T_1452_0 <= 1'h0;
    end else begin
      _T_1452_0 <= _T_95;
    end
    if (reset) begin
      _T_1452_1 <= 1'h0;
    end else begin
      _T_1452_1 <= _T_1452_0;
    end
    if (reset) begin
      _T_1452_2 <= 1'h0;
    end else begin
      _T_1452_2 <= _T_1452_1;
    end
    if (reset) begin
      _T_1452_3 <= 1'h0;
    end else begin
      _T_1452_3 <= _T_1452_2;
    end
    if (reset) begin
      _T_1462_0 <= 1'h0;
    end else begin
      _T_1462_0 <= _T_105;
    end
    if (reset) begin
      _T_1462_1 <= 1'h0;
    end else begin
      _T_1462_1 <= _T_1462_0;
    end
    if (reset) begin
      _T_1462_2 <= 1'h0;
    end else begin
      _T_1462_2 <= _T_1462_1;
    end
    if (reset) begin
      _T_1462_3 <= 1'h0;
    end else begin
      _T_1462_3 <= _T_1462_2;
    end
    if (reset) begin
      _T_1472_0 <= 1'h0;
    end else begin
      _T_1472_0 <= _T_115;
    end
    if (reset) begin
      _T_1472_1 <= 1'h0;
    end else begin
      _T_1472_1 <= _T_1472_0;
    end
    if (reset) begin
      _T_1472_2 <= 1'h0;
    end else begin
      _T_1472_2 <= _T_1472_1;
    end
    if (reset) begin
      _T_1472_3 <= 1'h0;
    end else begin
      _T_1472_3 <= _T_1472_2;
    end
    if (reset) begin
      _T_1482_0 <= 1'h0;
    end else begin
      _T_1482_0 <= _T_125;
    end
    if (reset) begin
      _T_1482_1 <= 1'h0;
    end else begin
      _T_1482_1 <= _T_1482_0;
    end
    if (reset) begin
      _T_1482_2 <= 1'h0;
    end else begin
      _T_1482_2 <= _T_1482_1;
    end
    if (reset) begin
      _T_1482_3 <= 1'h0;
    end else begin
      _T_1482_3 <= _T_1482_2;
    end
    if (reset) begin
      _T_1492_0 <= 1'h0;
    end else begin
      _T_1492_0 <= _T_135;
    end
    if (reset) begin
      _T_1492_1 <= 1'h0;
    end else begin
      _T_1492_1 <= _T_1492_0;
    end
    if (reset) begin
      _T_1492_2 <= 1'h0;
    end else begin
      _T_1492_2 <= _T_1492_1;
    end
    if (reset) begin
      _T_1492_3 <= 1'h0;
    end else begin
      _T_1492_3 <= _T_1492_2;
    end
    if (reset) begin
      _T_1502_0 <= 1'h0;
    end else begin
      _T_1502_0 <= _T_145;
    end
    if (reset) begin
      _T_1502_1 <= 1'h0;
    end else begin
      _T_1502_1 <= _T_1502_0;
    end
    if (reset) begin
      _T_1502_2 <= 1'h0;
    end else begin
      _T_1502_2 <= _T_1502_1;
    end
    if (reset) begin
      _T_1502_3 <= 1'h0;
    end else begin
      _T_1502_3 <= _T_1502_2;
    end
    if (reset) begin
      _T_1512_0 <= 1'h0;
    end else begin
      _T_1512_0 <= _T_155;
    end
    if (reset) begin
      _T_1512_1 <= 1'h0;
    end else begin
      _T_1512_1 <= _T_1512_0;
    end
    if (reset) begin
      _T_1512_2 <= 1'h0;
    end else begin
      _T_1512_2 <= _T_1512_1;
    end
    if (reset) begin
      _T_1512_3 <= 1'h0;
    end else begin
      _T_1512_3 <= _T_1512_2;
    end
    if (reset) begin
      _T_1522_0 <= 1'h0;
    end else begin
      _T_1522_0 <= _T_315;
    end
    if (reset) begin
      _T_1522_1 <= 1'h0;
    end else begin
      _T_1522_1 <= _T_1522_0;
    end
    if (reset) begin
      _T_1522_2 <= 1'h0;
    end else begin
      _T_1522_2 <= _T_1522_1;
    end
    if (reset) begin
      _T_1522_3 <= 1'h0;
    end else begin
      _T_1522_3 <= _T_1522_2;
    end
    if (reset) begin
      _T_1532_0 <= 1'h0;
    end else begin
      _T_1532_0 <= _T_475;
    end
    if (reset) begin
      _T_1532_1 <= 1'h0;
    end else begin
      _T_1532_1 <= _T_1532_0;
    end
    if (reset) begin
      _T_1532_2 <= 1'h0;
    end else begin
      _T_1532_2 <= _T_1532_1;
    end
    if (reset) begin
      _T_1532_3 <= 1'h0;
    end else begin
      _T_1532_3 <= _T_1532_2;
    end
    if (reset) begin
      _T_1542_0 <= 1'h0;
    end else begin
      _T_1542_0 <= _T_635;
    end
    if (reset) begin
      _T_1542_1 <= 1'h0;
    end else begin
      _T_1542_1 <= _T_1542_0;
    end
    if (reset) begin
      _T_1542_2 <= 1'h0;
    end else begin
      _T_1542_2 <= _T_1542_1;
    end
    if (reset) begin
      _T_1542_3 <= 1'h0;
    end else begin
      _T_1542_3 <= _T_1542_2;
    end
    if (reset) begin
      _T_1552_0 <= 1'h0;
    end else begin
      _T_1552_0 <= _T_795;
    end
    if (reset) begin
      _T_1552_1 <= 1'h0;
    end else begin
      _T_1552_1 <= _T_1552_0;
    end
    if (reset) begin
      _T_1552_2 <= 1'h0;
    end else begin
      _T_1552_2 <= _T_1552_1;
    end
    if (reset) begin
      _T_1552_3 <= 1'h0;
    end else begin
      _T_1552_3 <= _T_1552_2;
    end
    if (reset) begin
      _T_1562_0 <= 1'h0;
    end else begin
      _T_1562_0 <= _T_955;
    end
    if (reset) begin
      _T_1562_1 <= 1'h0;
    end else begin
      _T_1562_1 <= _T_1562_0;
    end
    if (reset) begin
      _T_1562_2 <= 1'h0;
    end else begin
      _T_1562_2 <= _T_1562_1;
    end
    if (reset) begin
      _T_1562_3 <= 1'h0;
    end else begin
      _T_1562_3 <= _T_1562_2;
    end
    if (reset) begin
      _T_1572_0 <= 1'h0;
    end else begin
      _T_1572_0 <= _T_1115;
    end
    if (reset) begin
      _T_1572_1 <= 1'h0;
    end else begin
      _T_1572_1 <= _T_1572_0;
    end
    if (reset) begin
      _T_1572_2 <= 1'h0;
    end else begin
      _T_1572_2 <= _T_1572_1;
    end
    if (reset) begin
      _T_1572_3 <= 1'h0;
    end else begin
      _T_1572_3 <= _T_1572_2;
    end
    if (reset) begin
      _T_1582_0 <= 1'h0;
    end else begin
      _T_1582_0 <= _T_1275;
    end
    if (reset) begin
      _T_1582_1 <= 1'h0;
    end else begin
      _T_1582_1 <= _T_1582_0;
    end
    if (reset) begin
      _T_1582_2 <= 1'h0;
    end else begin
      _T_1582_2 <= _T_1582_1;
    end
    if (reset) begin
      _T_1582_3 <= 1'h0;
    end else begin
      _T_1582_3 <= _T_1582_2;
    end
    if (reset) begin
      _T_1592_0 <= 1'h0;
    end else begin
      _T_1592_0 <= _T_1435;
    end
    if (reset) begin
      _T_1592_1 <= 1'h0;
    end else begin
      _T_1592_1 <= _T_1592_0;
    end
    if (reset) begin
      _T_1592_2 <= 1'h0;
    end else begin
      _T_1592_2 <= _T_1592_1;
    end
    if (reset) begin
      _T_1592_3 <= 1'h0;
    end else begin
      _T_1592_3 <= _T_1592_2;
    end
    if (reset) begin
      _T_1602_0 <= 1'h0;
    end else begin
      _T_1602_0 <= _T_1595;
    end
    if (reset) begin
      _T_1602_1 <= 1'h0;
    end else begin
      _T_1602_1 <= _T_1602_0;
    end
    if (reset) begin
      _T_1602_2 <= 1'h0;
    end else begin
      _T_1602_2 <= _T_1602_1;
    end
    if (reset) begin
      _T_1602_3 <= 1'h0;
    end else begin
      _T_1602_3 <= _T_1602_2;
    end
    if (reset) begin
      _T_1612_0 <= 1'h0;
    end else begin
      _T_1612_0 <= _T_105;
    end
    if (reset) begin
      _T_1612_1 <= 1'h0;
    end else begin
      _T_1612_1 <= _T_1612_0;
    end
    if (reset) begin
      _T_1612_2 <= 1'h0;
    end else begin
      _T_1612_2 <= _T_1612_1;
    end
    if (reset) begin
      _T_1612_3 <= 1'h0;
    end else begin
      _T_1612_3 <= _T_1612_2;
    end
    if (reset) begin
      _T_1622_0 <= 1'h0;
    end else begin
      _T_1622_0 <= _T_115;
    end
    if (reset) begin
      _T_1622_1 <= 1'h0;
    end else begin
      _T_1622_1 <= _T_1622_0;
    end
    if (reset) begin
      _T_1622_2 <= 1'h0;
    end else begin
      _T_1622_2 <= _T_1622_1;
    end
    if (reset) begin
      _T_1622_3 <= 1'h0;
    end else begin
      _T_1622_3 <= _T_1622_2;
    end
    if (reset) begin
      _T_1632_0 <= 1'h0;
    end else begin
      _T_1632_0 <= _T_125;
    end
    if (reset) begin
      _T_1632_1 <= 1'h0;
    end else begin
      _T_1632_1 <= _T_1632_0;
    end
    if (reset) begin
      _T_1632_2 <= 1'h0;
    end else begin
      _T_1632_2 <= _T_1632_1;
    end
    if (reset) begin
      _T_1632_3 <= 1'h0;
    end else begin
      _T_1632_3 <= _T_1632_2;
    end
    if (reset) begin
      _T_1642_0 <= 1'h0;
    end else begin
      _T_1642_0 <= _T_135;
    end
    if (reset) begin
      _T_1642_1 <= 1'h0;
    end else begin
      _T_1642_1 <= _T_1642_0;
    end
    if (reset) begin
      _T_1642_2 <= 1'h0;
    end else begin
      _T_1642_2 <= _T_1642_1;
    end
    if (reset) begin
      _T_1642_3 <= 1'h0;
    end else begin
      _T_1642_3 <= _T_1642_2;
    end
    if (reset) begin
      _T_1652_0 <= 1'h0;
    end else begin
      _T_1652_0 <= _T_145;
    end
    if (reset) begin
      _T_1652_1 <= 1'h0;
    end else begin
      _T_1652_1 <= _T_1652_0;
    end
    if (reset) begin
      _T_1652_2 <= 1'h0;
    end else begin
      _T_1652_2 <= _T_1652_1;
    end
    if (reset) begin
      _T_1652_3 <= 1'h0;
    end else begin
      _T_1652_3 <= _T_1652_2;
    end
    if (reset) begin
      _T_1662_0 <= 1'h0;
    end else begin
      _T_1662_0 <= _T_155;
    end
    if (reset) begin
      _T_1662_1 <= 1'h0;
    end else begin
      _T_1662_1 <= _T_1662_0;
    end
    if (reset) begin
      _T_1662_2 <= 1'h0;
    end else begin
      _T_1662_2 <= _T_1662_1;
    end
    if (reset) begin
      _T_1662_3 <= 1'h0;
    end else begin
      _T_1662_3 <= _T_1662_2;
    end
    if (reset) begin
      _T_1672_0 <= 1'h0;
    end else begin
      _T_1672_0 <= _T_315;
    end
    if (reset) begin
      _T_1672_1 <= 1'h0;
    end else begin
      _T_1672_1 <= _T_1672_0;
    end
    if (reset) begin
      _T_1672_2 <= 1'h0;
    end else begin
      _T_1672_2 <= _T_1672_1;
    end
    if (reset) begin
      _T_1672_3 <= 1'h0;
    end else begin
      _T_1672_3 <= _T_1672_2;
    end
    if (reset) begin
      _T_1682_0 <= 1'h0;
    end else begin
      _T_1682_0 <= _T_475;
    end
    if (reset) begin
      _T_1682_1 <= 1'h0;
    end else begin
      _T_1682_1 <= _T_1682_0;
    end
    if (reset) begin
      _T_1682_2 <= 1'h0;
    end else begin
      _T_1682_2 <= _T_1682_1;
    end
    if (reset) begin
      _T_1682_3 <= 1'h0;
    end else begin
      _T_1682_3 <= _T_1682_2;
    end
    if (reset) begin
      _T_1692_0 <= 1'h0;
    end else begin
      _T_1692_0 <= _T_635;
    end
    if (reset) begin
      _T_1692_1 <= 1'h0;
    end else begin
      _T_1692_1 <= _T_1692_0;
    end
    if (reset) begin
      _T_1692_2 <= 1'h0;
    end else begin
      _T_1692_2 <= _T_1692_1;
    end
    if (reset) begin
      _T_1692_3 <= 1'h0;
    end else begin
      _T_1692_3 <= _T_1692_2;
    end
    if (reset) begin
      _T_1702_0 <= 1'h0;
    end else begin
      _T_1702_0 <= _T_795;
    end
    if (reset) begin
      _T_1702_1 <= 1'h0;
    end else begin
      _T_1702_1 <= _T_1702_0;
    end
    if (reset) begin
      _T_1702_2 <= 1'h0;
    end else begin
      _T_1702_2 <= _T_1702_1;
    end
    if (reset) begin
      _T_1702_3 <= 1'h0;
    end else begin
      _T_1702_3 <= _T_1702_2;
    end
    if (reset) begin
      _T_1712_0 <= 1'h0;
    end else begin
      _T_1712_0 <= _T_955;
    end
    if (reset) begin
      _T_1712_1 <= 1'h0;
    end else begin
      _T_1712_1 <= _T_1712_0;
    end
    if (reset) begin
      _T_1712_2 <= 1'h0;
    end else begin
      _T_1712_2 <= _T_1712_1;
    end
    if (reset) begin
      _T_1712_3 <= 1'h0;
    end else begin
      _T_1712_3 <= _T_1712_2;
    end
    if (reset) begin
      _T_1722_0 <= 1'h0;
    end else begin
      _T_1722_0 <= _T_1115;
    end
    if (reset) begin
      _T_1722_1 <= 1'h0;
    end else begin
      _T_1722_1 <= _T_1722_0;
    end
    if (reset) begin
      _T_1722_2 <= 1'h0;
    end else begin
      _T_1722_2 <= _T_1722_1;
    end
    if (reset) begin
      _T_1722_3 <= 1'h0;
    end else begin
      _T_1722_3 <= _T_1722_2;
    end
    if (reset) begin
      _T_1732_0 <= 1'h0;
    end else begin
      _T_1732_0 <= _T_1275;
    end
    if (reset) begin
      _T_1732_1 <= 1'h0;
    end else begin
      _T_1732_1 <= _T_1732_0;
    end
    if (reset) begin
      _T_1732_2 <= 1'h0;
    end else begin
      _T_1732_2 <= _T_1732_1;
    end
    if (reset) begin
      _T_1732_3 <= 1'h0;
    end else begin
      _T_1732_3 <= _T_1732_2;
    end
    if (reset) begin
      _T_1742_0 <= 1'h0;
    end else begin
      _T_1742_0 <= _T_1435;
    end
    if (reset) begin
      _T_1742_1 <= 1'h0;
    end else begin
      _T_1742_1 <= _T_1742_0;
    end
    if (reset) begin
      _T_1742_2 <= 1'h0;
    end else begin
      _T_1742_2 <= _T_1742_1;
    end
    if (reset) begin
      _T_1742_3 <= 1'h0;
    end else begin
      _T_1742_3 <= _T_1742_2;
    end
    if (reset) begin
      _T_1752_0 <= 1'h0;
    end else begin
      _T_1752_0 <= _T_1595;
    end
    if (reset) begin
      _T_1752_1 <= 1'h0;
    end else begin
      _T_1752_1 <= _T_1752_0;
    end
    if (reset) begin
      _T_1752_2 <= 1'h0;
    end else begin
      _T_1752_2 <= _T_1752_1;
    end
    if (reset) begin
      _T_1752_3 <= 1'h0;
    end else begin
      _T_1752_3 <= _T_1752_2;
    end
    if (reset) begin
      _T_1762_0 <= 1'h0;
    end else begin
      _T_1762_0 <= _T_1755;
    end
    if (reset) begin
      _T_1762_1 <= 1'h0;
    end else begin
      _T_1762_1 <= _T_1762_0;
    end
    if (reset) begin
      _T_1762_2 <= 1'h0;
    end else begin
      _T_1762_2 <= _T_1762_1;
    end
    if (reset) begin
      _T_1762_3 <= 1'h0;
    end else begin
      _T_1762_3 <= _T_1762_2;
    end
    if (reset) begin
      _T_1772_0 <= 1'h0;
    end else begin
      _T_1772_0 <= _T_115;
    end
    if (reset) begin
      _T_1772_1 <= 1'h0;
    end else begin
      _T_1772_1 <= _T_1772_0;
    end
    if (reset) begin
      _T_1772_2 <= 1'h0;
    end else begin
      _T_1772_2 <= _T_1772_1;
    end
    if (reset) begin
      _T_1772_3 <= 1'h0;
    end else begin
      _T_1772_3 <= _T_1772_2;
    end
    if (reset) begin
      _T_1782_0 <= 1'h0;
    end else begin
      _T_1782_0 <= _T_125;
    end
    if (reset) begin
      _T_1782_1 <= 1'h0;
    end else begin
      _T_1782_1 <= _T_1782_0;
    end
    if (reset) begin
      _T_1782_2 <= 1'h0;
    end else begin
      _T_1782_2 <= _T_1782_1;
    end
    if (reset) begin
      _T_1782_3 <= 1'h0;
    end else begin
      _T_1782_3 <= _T_1782_2;
    end
    if (reset) begin
      _T_1792_0 <= 1'h0;
    end else begin
      _T_1792_0 <= _T_135;
    end
    if (reset) begin
      _T_1792_1 <= 1'h0;
    end else begin
      _T_1792_1 <= _T_1792_0;
    end
    if (reset) begin
      _T_1792_2 <= 1'h0;
    end else begin
      _T_1792_2 <= _T_1792_1;
    end
    if (reset) begin
      _T_1792_3 <= 1'h0;
    end else begin
      _T_1792_3 <= _T_1792_2;
    end
    if (reset) begin
      _T_1802_0 <= 1'h0;
    end else begin
      _T_1802_0 <= _T_145;
    end
    if (reset) begin
      _T_1802_1 <= 1'h0;
    end else begin
      _T_1802_1 <= _T_1802_0;
    end
    if (reset) begin
      _T_1802_2 <= 1'h0;
    end else begin
      _T_1802_2 <= _T_1802_1;
    end
    if (reset) begin
      _T_1802_3 <= 1'h0;
    end else begin
      _T_1802_3 <= _T_1802_2;
    end
    if (reset) begin
      _T_1812_0 <= 1'h0;
    end else begin
      _T_1812_0 <= _T_155;
    end
    if (reset) begin
      _T_1812_1 <= 1'h0;
    end else begin
      _T_1812_1 <= _T_1812_0;
    end
    if (reset) begin
      _T_1812_2 <= 1'h0;
    end else begin
      _T_1812_2 <= _T_1812_1;
    end
    if (reset) begin
      _T_1812_3 <= 1'h0;
    end else begin
      _T_1812_3 <= _T_1812_2;
    end
    if (reset) begin
      _T_1822_0 <= 1'h0;
    end else begin
      _T_1822_0 <= _T_315;
    end
    if (reset) begin
      _T_1822_1 <= 1'h0;
    end else begin
      _T_1822_1 <= _T_1822_0;
    end
    if (reset) begin
      _T_1822_2 <= 1'h0;
    end else begin
      _T_1822_2 <= _T_1822_1;
    end
    if (reset) begin
      _T_1822_3 <= 1'h0;
    end else begin
      _T_1822_3 <= _T_1822_2;
    end
    if (reset) begin
      _T_1832_0 <= 1'h0;
    end else begin
      _T_1832_0 <= _T_475;
    end
    if (reset) begin
      _T_1832_1 <= 1'h0;
    end else begin
      _T_1832_1 <= _T_1832_0;
    end
    if (reset) begin
      _T_1832_2 <= 1'h0;
    end else begin
      _T_1832_2 <= _T_1832_1;
    end
    if (reset) begin
      _T_1832_3 <= 1'h0;
    end else begin
      _T_1832_3 <= _T_1832_2;
    end
    if (reset) begin
      _T_1842_0 <= 1'h0;
    end else begin
      _T_1842_0 <= _T_635;
    end
    if (reset) begin
      _T_1842_1 <= 1'h0;
    end else begin
      _T_1842_1 <= _T_1842_0;
    end
    if (reset) begin
      _T_1842_2 <= 1'h0;
    end else begin
      _T_1842_2 <= _T_1842_1;
    end
    if (reset) begin
      _T_1842_3 <= 1'h0;
    end else begin
      _T_1842_3 <= _T_1842_2;
    end
    if (reset) begin
      _T_1852_0 <= 1'h0;
    end else begin
      _T_1852_0 <= _T_795;
    end
    if (reset) begin
      _T_1852_1 <= 1'h0;
    end else begin
      _T_1852_1 <= _T_1852_0;
    end
    if (reset) begin
      _T_1852_2 <= 1'h0;
    end else begin
      _T_1852_2 <= _T_1852_1;
    end
    if (reset) begin
      _T_1852_3 <= 1'h0;
    end else begin
      _T_1852_3 <= _T_1852_2;
    end
    if (reset) begin
      _T_1862_0 <= 1'h0;
    end else begin
      _T_1862_0 <= _T_955;
    end
    if (reset) begin
      _T_1862_1 <= 1'h0;
    end else begin
      _T_1862_1 <= _T_1862_0;
    end
    if (reset) begin
      _T_1862_2 <= 1'h0;
    end else begin
      _T_1862_2 <= _T_1862_1;
    end
    if (reset) begin
      _T_1862_3 <= 1'h0;
    end else begin
      _T_1862_3 <= _T_1862_2;
    end
    if (reset) begin
      _T_1872_0 <= 1'h0;
    end else begin
      _T_1872_0 <= _T_1115;
    end
    if (reset) begin
      _T_1872_1 <= 1'h0;
    end else begin
      _T_1872_1 <= _T_1872_0;
    end
    if (reset) begin
      _T_1872_2 <= 1'h0;
    end else begin
      _T_1872_2 <= _T_1872_1;
    end
    if (reset) begin
      _T_1872_3 <= 1'h0;
    end else begin
      _T_1872_3 <= _T_1872_2;
    end
    if (reset) begin
      _T_1882_0 <= 1'h0;
    end else begin
      _T_1882_0 <= _T_1275;
    end
    if (reset) begin
      _T_1882_1 <= 1'h0;
    end else begin
      _T_1882_1 <= _T_1882_0;
    end
    if (reset) begin
      _T_1882_2 <= 1'h0;
    end else begin
      _T_1882_2 <= _T_1882_1;
    end
    if (reset) begin
      _T_1882_3 <= 1'h0;
    end else begin
      _T_1882_3 <= _T_1882_2;
    end
    if (reset) begin
      _T_1892_0 <= 1'h0;
    end else begin
      _T_1892_0 <= _T_1435;
    end
    if (reset) begin
      _T_1892_1 <= 1'h0;
    end else begin
      _T_1892_1 <= _T_1892_0;
    end
    if (reset) begin
      _T_1892_2 <= 1'h0;
    end else begin
      _T_1892_2 <= _T_1892_1;
    end
    if (reset) begin
      _T_1892_3 <= 1'h0;
    end else begin
      _T_1892_3 <= _T_1892_2;
    end
    if (reset) begin
      _T_1902_0 <= 1'h0;
    end else begin
      _T_1902_0 <= _T_1595;
    end
    if (reset) begin
      _T_1902_1 <= 1'h0;
    end else begin
      _T_1902_1 <= _T_1902_0;
    end
    if (reset) begin
      _T_1902_2 <= 1'h0;
    end else begin
      _T_1902_2 <= _T_1902_1;
    end
    if (reset) begin
      _T_1902_3 <= 1'h0;
    end else begin
      _T_1902_3 <= _T_1902_2;
    end
    if (reset) begin
      _T_1912_0 <= 1'h0;
    end else begin
      _T_1912_0 <= _T_1755;
    end
    if (reset) begin
      _T_1912_1 <= 1'h0;
    end else begin
      _T_1912_1 <= _T_1912_0;
    end
    if (reset) begin
      _T_1912_2 <= 1'h0;
    end else begin
      _T_1912_2 <= _T_1912_1;
    end
    if (reset) begin
      _T_1912_3 <= 1'h0;
    end else begin
      _T_1912_3 <= _T_1912_2;
    end
    if (reset) begin
      _T_1922_0 <= 1'h0;
    end else begin
      _T_1922_0 <= _T_1915;
    end
    if (reset) begin
      _T_1922_1 <= 1'h0;
    end else begin
      _T_1922_1 <= _T_1922_0;
    end
    if (reset) begin
      _T_1922_2 <= 1'h0;
    end else begin
      _T_1922_2 <= _T_1922_1;
    end
    if (reset) begin
      _T_1922_3 <= 1'h0;
    end else begin
      _T_1922_3 <= _T_1922_2;
    end
    if (reset) begin
      _T_1932_0 <= 1'h0;
    end else begin
      _T_1932_0 <= _T_125;
    end
    if (reset) begin
      _T_1932_1 <= 1'h0;
    end else begin
      _T_1932_1 <= _T_1932_0;
    end
    if (reset) begin
      _T_1932_2 <= 1'h0;
    end else begin
      _T_1932_2 <= _T_1932_1;
    end
    if (reset) begin
      _T_1932_3 <= 1'h0;
    end else begin
      _T_1932_3 <= _T_1932_2;
    end
    if (reset) begin
      _T_1942_0 <= 1'h0;
    end else begin
      _T_1942_0 <= _T_135;
    end
    if (reset) begin
      _T_1942_1 <= 1'h0;
    end else begin
      _T_1942_1 <= _T_1942_0;
    end
    if (reset) begin
      _T_1942_2 <= 1'h0;
    end else begin
      _T_1942_2 <= _T_1942_1;
    end
    if (reset) begin
      _T_1942_3 <= 1'h0;
    end else begin
      _T_1942_3 <= _T_1942_2;
    end
    if (reset) begin
      _T_1952_0 <= 1'h0;
    end else begin
      _T_1952_0 <= _T_145;
    end
    if (reset) begin
      _T_1952_1 <= 1'h0;
    end else begin
      _T_1952_1 <= _T_1952_0;
    end
    if (reset) begin
      _T_1952_2 <= 1'h0;
    end else begin
      _T_1952_2 <= _T_1952_1;
    end
    if (reset) begin
      _T_1952_3 <= 1'h0;
    end else begin
      _T_1952_3 <= _T_1952_2;
    end
    if (reset) begin
      _T_1962_0 <= 1'h0;
    end else begin
      _T_1962_0 <= _T_155;
    end
    if (reset) begin
      _T_1962_1 <= 1'h0;
    end else begin
      _T_1962_1 <= _T_1962_0;
    end
    if (reset) begin
      _T_1962_2 <= 1'h0;
    end else begin
      _T_1962_2 <= _T_1962_1;
    end
    if (reset) begin
      _T_1962_3 <= 1'h0;
    end else begin
      _T_1962_3 <= _T_1962_2;
    end
    if (reset) begin
      _T_1972_0 <= 1'h0;
    end else begin
      _T_1972_0 <= _T_315;
    end
    if (reset) begin
      _T_1972_1 <= 1'h0;
    end else begin
      _T_1972_1 <= _T_1972_0;
    end
    if (reset) begin
      _T_1972_2 <= 1'h0;
    end else begin
      _T_1972_2 <= _T_1972_1;
    end
    if (reset) begin
      _T_1972_3 <= 1'h0;
    end else begin
      _T_1972_3 <= _T_1972_2;
    end
    if (reset) begin
      _T_1982_0 <= 1'h0;
    end else begin
      _T_1982_0 <= _T_475;
    end
    if (reset) begin
      _T_1982_1 <= 1'h0;
    end else begin
      _T_1982_1 <= _T_1982_0;
    end
    if (reset) begin
      _T_1982_2 <= 1'h0;
    end else begin
      _T_1982_2 <= _T_1982_1;
    end
    if (reset) begin
      _T_1982_3 <= 1'h0;
    end else begin
      _T_1982_3 <= _T_1982_2;
    end
    if (reset) begin
      _T_1992_0 <= 1'h0;
    end else begin
      _T_1992_0 <= _T_635;
    end
    if (reset) begin
      _T_1992_1 <= 1'h0;
    end else begin
      _T_1992_1 <= _T_1992_0;
    end
    if (reset) begin
      _T_1992_2 <= 1'h0;
    end else begin
      _T_1992_2 <= _T_1992_1;
    end
    if (reset) begin
      _T_1992_3 <= 1'h0;
    end else begin
      _T_1992_3 <= _T_1992_2;
    end
    if (reset) begin
      _T_2002_0 <= 1'h0;
    end else begin
      _T_2002_0 <= _T_795;
    end
    if (reset) begin
      _T_2002_1 <= 1'h0;
    end else begin
      _T_2002_1 <= _T_2002_0;
    end
    if (reset) begin
      _T_2002_2 <= 1'h0;
    end else begin
      _T_2002_2 <= _T_2002_1;
    end
    if (reset) begin
      _T_2002_3 <= 1'h0;
    end else begin
      _T_2002_3 <= _T_2002_2;
    end
    if (reset) begin
      _T_2012_0 <= 1'h0;
    end else begin
      _T_2012_0 <= _T_955;
    end
    if (reset) begin
      _T_2012_1 <= 1'h0;
    end else begin
      _T_2012_1 <= _T_2012_0;
    end
    if (reset) begin
      _T_2012_2 <= 1'h0;
    end else begin
      _T_2012_2 <= _T_2012_1;
    end
    if (reset) begin
      _T_2012_3 <= 1'h0;
    end else begin
      _T_2012_3 <= _T_2012_2;
    end
    if (reset) begin
      _T_2022_0 <= 1'h0;
    end else begin
      _T_2022_0 <= _T_1115;
    end
    if (reset) begin
      _T_2022_1 <= 1'h0;
    end else begin
      _T_2022_1 <= _T_2022_0;
    end
    if (reset) begin
      _T_2022_2 <= 1'h0;
    end else begin
      _T_2022_2 <= _T_2022_1;
    end
    if (reset) begin
      _T_2022_3 <= 1'h0;
    end else begin
      _T_2022_3 <= _T_2022_2;
    end
    if (reset) begin
      _T_2032_0 <= 1'h0;
    end else begin
      _T_2032_0 <= _T_1275;
    end
    if (reset) begin
      _T_2032_1 <= 1'h0;
    end else begin
      _T_2032_1 <= _T_2032_0;
    end
    if (reset) begin
      _T_2032_2 <= 1'h0;
    end else begin
      _T_2032_2 <= _T_2032_1;
    end
    if (reset) begin
      _T_2032_3 <= 1'h0;
    end else begin
      _T_2032_3 <= _T_2032_2;
    end
    if (reset) begin
      _T_2042_0 <= 1'h0;
    end else begin
      _T_2042_0 <= _T_1435;
    end
    if (reset) begin
      _T_2042_1 <= 1'h0;
    end else begin
      _T_2042_1 <= _T_2042_0;
    end
    if (reset) begin
      _T_2042_2 <= 1'h0;
    end else begin
      _T_2042_2 <= _T_2042_1;
    end
    if (reset) begin
      _T_2042_3 <= 1'h0;
    end else begin
      _T_2042_3 <= _T_2042_2;
    end
    if (reset) begin
      _T_2052_0 <= 1'h0;
    end else begin
      _T_2052_0 <= _T_1595;
    end
    if (reset) begin
      _T_2052_1 <= 1'h0;
    end else begin
      _T_2052_1 <= _T_2052_0;
    end
    if (reset) begin
      _T_2052_2 <= 1'h0;
    end else begin
      _T_2052_2 <= _T_2052_1;
    end
    if (reset) begin
      _T_2052_3 <= 1'h0;
    end else begin
      _T_2052_3 <= _T_2052_2;
    end
    if (reset) begin
      _T_2062_0 <= 1'h0;
    end else begin
      _T_2062_0 <= _T_1755;
    end
    if (reset) begin
      _T_2062_1 <= 1'h0;
    end else begin
      _T_2062_1 <= _T_2062_0;
    end
    if (reset) begin
      _T_2062_2 <= 1'h0;
    end else begin
      _T_2062_2 <= _T_2062_1;
    end
    if (reset) begin
      _T_2062_3 <= 1'h0;
    end else begin
      _T_2062_3 <= _T_2062_2;
    end
    if (reset) begin
      _T_2072_0 <= 1'h0;
    end else begin
      _T_2072_0 <= _T_1915;
    end
    if (reset) begin
      _T_2072_1 <= 1'h0;
    end else begin
      _T_2072_1 <= _T_2072_0;
    end
    if (reset) begin
      _T_2072_2 <= 1'h0;
    end else begin
      _T_2072_2 <= _T_2072_1;
    end
    if (reset) begin
      _T_2072_3 <= 1'h0;
    end else begin
      _T_2072_3 <= _T_2072_2;
    end
    if (reset) begin
      _T_2082_0 <= 1'h0;
    end else begin
      _T_2082_0 <= _T_2075;
    end
    if (reset) begin
      _T_2082_1 <= 1'h0;
    end else begin
      _T_2082_1 <= _T_2082_0;
    end
    if (reset) begin
      _T_2082_2 <= 1'h0;
    end else begin
      _T_2082_2 <= _T_2082_1;
    end
    if (reset) begin
      _T_2082_3 <= 1'h0;
    end else begin
      _T_2082_3 <= _T_2082_2;
    end
    if (reset) begin
      _T_2092_0 <= 1'h0;
    end else begin
      _T_2092_0 <= _T_135;
    end
    if (reset) begin
      _T_2092_1 <= 1'h0;
    end else begin
      _T_2092_1 <= _T_2092_0;
    end
    if (reset) begin
      _T_2092_2 <= 1'h0;
    end else begin
      _T_2092_2 <= _T_2092_1;
    end
    if (reset) begin
      _T_2092_3 <= 1'h0;
    end else begin
      _T_2092_3 <= _T_2092_2;
    end
    if (reset) begin
      _T_2102_0 <= 1'h0;
    end else begin
      _T_2102_0 <= _T_145;
    end
    if (reset) begin
      _T_2102_1 <= 1'h0;
    end else begin
      _T_2102_1 <= _T_2102_0;
    end
    if (reset) begin
      _T_2102_2 <= 1'h0;
    end else begin
      _T_2102_2 <= _T_2102_1;
    end
    if (reset) begin
      _T_2102_3 <= 1'h0;
    end else begin
      _T_2102_3 <= _T_2102_2;
    end
    if (reset) begin
      _T_2112_0 <= 1'h0;
    end else begin
      _T_2112_0 <= _T_155;
    end
    if (reset) begin
      _T_2112_1 <= 1'h0;
    end else begin
      _T_2112_1 <= _T_2112_0;
    end
    if (reset) begin
      _T_2112_2 <= 1'h0;
    end else begin
      _T_2112_2 <= _T_2112_1;
    end
    if (reset) begin
      _T_2112_3 <= 1'h0;
    end else begin
      _T_2112_3 <= _T_2112_2;
    end
    if (reset) begin
      _T_2122_0 <= 1'h0;
    end else begin
      _T_2122_0 <= _T_315;
    end
    if (reset) begin
      _T_2122_1 <= 1'h0;
    end else begin
      _T_2122_1 <= _T_2122_0;
    end
    if (reset) begin
      _T_2122_2 <= 1'h0;
    end else begin
      _T_2122_2 <= _T_2122_1;
    end
    if (reset) begin
      _T_2122_3 <= 1'h0;
    end else begin
      _T_2122_3 <= _T_2122_2;
    end
    if (reset) begin
      _T_2132_0 <= 1'h0;
    end else begin
      _T_2132_0 <= _T_475;
    end
    if (reset) begin
      _T_2132_1 <= 1'h0;
    end else begin
      _T_2132_1 <= _T_2132_0;
    end
    if (reset) begin
      _T_2132_2 <= 1'h0;
    end else begin
      _T_2132_2 <= _T_2132_1;
    end
    if (reset) begin
      _T_2132_3 <= 1'h0;
    end else begin
      _T_2132_3 <= _T_2132_2;
    end
    if (reset) begin
      _T_2142_0 <= 1'h0;
    end else begin
      _T_2142_0 <= _T_635;
    end
    if (reset) begin
      _T_2142_1 <= 1'h0;
    end else begin
      _T_2142_1 <= _T_2142_0;
    end
    if (reset) begin
      _T_2142_2 <= 1'h0;
    end else begin
      _T_2142_2 <= _T_2142_1;
    end
    if (reset) begin
      _T_2142_3 <= 1'h0;
    end else begin
      _T_2142_3 <= _T_2142_2;
    end
    if (reset) begin
      _T_2152_0 <= 1'h0;
    end else begin
      _T_2152_0 <= _T_795;
    end
    if (reset) begin
      _T_2152_1 <= 1'h0;
    end else begin
      _T_2152_1 <= _T_2152_0;
    end
    if (reset) begin
      _T_2152_2 <= 1'h0;
    end else begin
      _T_2152_2 <= _T_2152_1;
    end
    if (reset) begin
      _T_2152_3 <= 1'h0;
    end else begin
      _T_2152_3 <= _T_2152_2;
    end
    if (reset) begin
      _T_2162_0 <= 1'h0;
    end else begin
      _T_2162_0 <= _T_955;
    end
    if (reset) begin
      _T_2162_1 <= 1'h0;
    end else begin
      _T_2162_1 <= _T_2162_0;
    end
    if (reset) begin
      _T_2162_2 <= 1'h0;
    end else begin
      _T_2162_2 <= _T_2162_1;
    end
    if (reset) begin
      _T_2162_3 <= 1'h0;
    end else begin
      _T_2162_3 <= _T_2162_2;
    end
    if (reset) begin
      _T_2172_0 <= 1'h0;
    end else begin
      _T_2172_0 <= _T_1115;
    end
    if (reset) begin
      _T_2172_1 <= 1'h0;
    end else begin
      _T_2172_1 <= _T_2172_0;
    end
    if (reset) begin
      _T_2172_2 <= 1'h0;
    end else begin
      _T_2172_2 <= _T_2172_1;
    end
    if (reset) begin
      _T_2172_3 <= 1'h0;
    end else begin
      _T_2172_3 <= _T_2172_2;
    end
    if (reset) begin
      _T_2182_0 <= 1'h0;
    end else begin
      _T_2182_0 <= _T_1275;
    end
    if (reset) begin
      _T_2182_1 <= 1'h0;
    end else begin
      _T_2182_1 <= _T_2182_0;
    end
    if (reset) begin
      _T_2182_2 <= 1'h0;
    end else begin
      _T_2182_2 <= _T_2182_1;
    end
    if (reset) begin
      _T_2182_3 <= 1'h0;
    end else begin
      _T_2182_3 <= _T_2182_2;
    end
    if (reset) begin
      _T_2192_0 <= 1'h0;
    end else begin
      _T_2192_0 <= _T_1435;
    end
    if (reset) begin
      _T_2192_1 <= 1'h0;
    end else begin
      _T_2192_1 <= _T_2192_0;
    end
    if (reset) begin
      _T_2192_2 <= 1'h0;
    end else begin
      _T_2192_2 <= _T_2192_1;
    end
    if (reset) begin
      _T_2192_3 <= 1'h0;
    end else begin
      _T_2192_3 <= _T_2192_2;
    end
    if (reset) begin
      _T_2202_0 <= 1'h0;
    end else begin
      _T_2202_0 <= _T_1595;
    end
    if (reset) begin
      _T_2202_1 <= 1'h0;
    end else begin
      _T_2202_1 <= _T_2202_0;
    end
    if (reset) begin
      _T_2202_2 <= 1'h0;
    end else begin
      _T_2202_2 <= _T_2202_1;
    end
    if (reset) begin
      _T_2202_3 <= 1'h0;
    end else begin
      _T_2202_3 <= _T_2202_2;
    end
    if (reset) begin
      _T_2212_0 <= 1'h0;
    end else begin
      _T_2212_0 <= _T_1755;
    end
    if (reset) begin
      _T_2212_1 <= 1'h0;
    end else begin
      _T_2212_1 <= _T_2212_0;
    end
    if (reset) begin
      _T_2212_2 <= 1'h0;
    end else begin
      _T_2212_2 <= _T_2212_1;
    end
    if (reset) begin
      _T_2212_3 <= 1'h0;
    end else begin
      _T_2212_3 <= _T_2212_2;
    end
    if (reset) begin
      _T_2222_0 <= 1'h0;
    end else begin
      _T_2222_0 <= _T_1915;
    end
    if (reset) begin
      _T_2222_1 <= 1'h0;
    end else begin
      _T_2222_1 <= _T_2222_0;
    end
    if (reset) begin
      _T_2222_2 <= 1'h0;
    end else begin
      _T_2222_2 <= _T_2222_1;
    end
    if (reset) begin
      _T_2222_3 <= 1'h0;
    end else begin
      _T_2222_3 <= _T_2222_2;
    end
    if (reset) begin
      _T_2232_0 <= 1'h0;
    end else begin
      _T_2232_0 <= _T_2075;
    end
    if (reset) begin
      _T_2232_1 <= 1'h0;
    end else begin
      _T_2232_1 <= _T_2232_0;
    end
    if (reset) begin
      _T_2232_2 <= 1'h0;
    end else begin
      _T_2232_2 <= _T_2232_1;
    end
    if (reset) begin
      _T_2232_3 <= 1'h0;
    end else begin
      _T_2232_3 <= _T_2232_2;
    end
    if (reset) begin
      _T_2242_0 <= 1'h0;
    end else begin
      _T_2242_0 <= _T_2235;
    end
    if (reset) begin
      _T_2242_1 <= 1'h0;
    end else begin
      _T_2242_1 <= _T_2242_0;
    end
    if (reset) begin
      _T_2242_2 <= 1'h0;
    end else begin
      _T_2242_2 <= _T_2242_1;
    end
    if (reset) begin
      _T_2242_3 <= 1'h0;
    end else begin
      _T_2242_3 <= _T_2242_2;
    end
    if (reset) begin
      _T_2252_0 <= 1'h0;
    end else begin
      _T_2252_0 <= _T_145;
    end
    if (reset) begin
      _T_2252_1 <= 1'h0;
    end else begin
      _T_2252_1 <= _T_2252_0;
    end
    if (reset) begin
      _T_2252_2 <= 1'h0;
    end else begin
      _T_2252_2 <= _T_2252_1;
    end
    if (reset) begin
      _T_2252_3 <= 1'h0;
    end else begin
      _T_2252_3 <= _T_2252_2;
    end
    if (reset) begin
      _T_2262_0 <= 1'h0;
    end else begin
      _T_2262_0 <= _T_155;
    end
    if (reset) begin
      _T_2262_1 <= 1'h0;
    end else begin
      _T_2262_1 <= _T_2262_0;
    end
    if (reset) begin
      _T_2262_2 <= 1'h0;
    end else begin
      _T_2262_2 <= _T_2262_1;
    end
    if (reset) begin
      _T_2262_3 <= 1'h0;
    end else begin
      _T_2262_3 <= _T_2262_2;
    end
    if (reset) begin
      _T_2272_0 <= 1'h0;
    end else begin
      _T_2272_0 <= _T_315;
    end
    if (reset) begin
      _T_2272_1 <= 1'h0;
    end else begin
      _T_2272_1 <= _T_2272_0;
    end
    if (reset) begin
      _T_2272_2 <= 1'h0;
    end else begin
      _T_2272_2 <= _T_2272_1;
    end
    if (reset) begin
      _T_2272_3 <= 1'h0;
    end else begin
      _T_2272_3 <= _T_2272_2;
    end
    if (reset) begin
      _T_2282_0 <= 1'h0;
    end else begin
      _T_2282_0 <= _T_475;
    end
    if (reset) begin
      _T_2282_1 <= 1'h0;
    end else begin
      _T_2282_1 <= _T_2282_0;
    end
    if (reset) begin
      _T_2282_2 <= 1'h0;
    end else begin
      _T_2282_2 <= _T_2282_1;
    end
    if (reset) begin
      _T_2282_3 <= 1'h0;
    end else begin
      _T_2282_3 <= _T_2282_2;
    end
    if (reset) begin
      _T_2292_0 <= 1'h0;
    end else begin
      _T_2292_0 <= _T_635;
    end
    if (reset) begin
      _T_2292_1 <= 1'h0;
    end else begin
      _T_2292_1 <= _T_2292_0;
    end
    if (reset) begin
      _T_2292_2 <= 1'h0;
    end else begin
      _T_2292_2 <= _T_2292_1;
    end
    if (reset) begin
      _T_2292_3 <= 1'h0;
    end else begin
      _T_2292_3 <= _T_2292_2;
    end
    if (reset) begin
      _T_2302_0 <= 1'h0;
    end else begin
      _T_2302_0 <= _T_795;
    end
    if (reset) begin
      _T_2302_1 <= 1'h0;
    end else begin
      _T_2302_1 <= _T_2302_0;
    end
    if (reset) begin
      _T_2302_2 <= 1'h0;
    end else begin
      _T_2302_2 <= _T_2302_1;
    end
    if (reset) begin
      _T_2302_3 <= 1'h0;
    end else begin
      _T_2302_3 <= _T_2302_2;
    end
    if (reset) begin
      _T_2312_0 <= 1'h0;
    end else begin
      _T_2312_0 <= _T_955;
    end
    if (reset) begin
      _T_2312_1 <= 1'h0;
    end else begin
      _T_2312_1 <= _T_2312_0;
    end
    if (reset) begin
      _T_2312_2 <= 1'h0;
    end else begin
      _T_2312_2 <= _T_2312_1;
    end
    if (reset) begin
      _T_2312_3 <= 1'h0;
    end else begin
      _T_2312_3 <= _T_2312_2;
    end
    if (reset) begin
      _T_2322_0 <= 1'h0;
    end else begin
      _T_2322_0 <= _T_1115;
    end
    if (reset) begin
      _T_2322_1 <= 1'h0;
    end else begin
      _T_2322_1 <= _T_2322_0;
    end
    if (reset) begin
      _T_2322_2 <= 1'h0;
    end else begin
      _T_2322_2 <= _T_2322_1;
    end
    if (reset) begin
      _T_2322_3 <= 1'h0;
    end else begin
      _T_2322_3 <= _T_2322_2;
    end
    if (reset) begin
      _T_2332_0 <= 1'h0;
    end else begin
      _T_2332_0 <= _T_1275;
    end
    if (reset) begin
      _T_2332_1 <= 1'h0;
    end else begin
      _T_2332_1 <= _T_2332_0;
    end
    if (reset) begin
      _T_2332_2 <= 1'h0;
    end else begin
      _T_2332_2 <= _T_2332_1;
    end
    if (reset) begin
      _T_2332_3 <= 1'h0;
    end else begin
      _T_2332_3 <= _T_2332_2;
    end
    if (reset) begin
      _T_2342_0 <= 1'h0;
    end else begin
      _T_2342_0 <= _T_1435;
    end
    if (reset) begin
      _T_2342_1 <= 1'h0;
    end else begin
      _T_2342_1 <= _T_2342_0;
    end
    if (reset) begin
      _T_2342_2 <= 1'h0;
    end else begin
      _T_2342_2 <= _T_2342_1;
    end
    if (reset) begin
      _T_2342_3 <= 1'h0;
    end else begin
      _T_2342_3 <= _T_2342_2;
    end
    if (reset) begin
      _T_2352_0 <= 1'h0;
    end else begin
      _T_2352_0 <= _T_1595;
    end
    if (reset) begin
      _T_2352_1 <= 1'h0;
    end else begin
      _T_2352_1 <= _T_2352_0;
    end
    if (reset) begin
      _T_2352_2 <= 1'h0;
    end else begin
      _T_2352_2 <= _T_2352_1;
    end
    if (reset) begin
      _T_2352_3 <= 1'h0;
    end else begin
      _T_2352_3 <= _T_2352_2;
    end
    if (reset) begin
      _T_2362_0 <= 1'h0;
    end else begin
      _T_2362_0 <= _T_1755;
    end
    if (reset) begin
      _T_2362_1 <= 1'h0;
    end else begin
      _T_2362_1 <= _T_2362_0;
    end
    if (reset) begin
      _T_2362_2 <= 1'h0;
    end else begin
      _T_2362_2 <= _T_2362_1;
    end
    if (reset) begin
      _T_2362_3 <= 1'h0;
    end else begin
      _T_2362_3 <= _T_2362_2;
    end
    if (reset) begin
      _T_2372_0 <= 1'h0;
    end else begin
      _T_2372_0 <= _T_1915;
    end
    if (reset) begin
      _T_2372_1 <= 1'h0;
    end else begin
      _T_2372_1 <= _T_2372_0;
    end
    if (reset) begin
      _T_2372_2 <= 1'h0;
    end else begin
      _T_2372_2 <= _T_2372_1;
    end
    if (reset) begin
      _T_2372_3 <= 1'h0;
    end else begin
      _T_2372_3 <= _T_2372_2;
    end
    if (reset) begin
      _T_2382_0 <= 1'h0;
    end else begin
      _T_2382_0 <= _T_2075;
    end
    if (reset) begin
      _T_2382_1 <= 1'h0;
    end else begin
      _T_2382_1 <= _T_2382_0;
    end
    if (reset) begin
      _T_2382_2 <= 1'h0;
    end else begin
      _T_2382_2 <= _T_2382_1;
    end
    if (reset) begin
      _T_2382_3 <= 1'h0;
    end else begin
      _T_2382_3 <= _T_2382_2;
    end
    if (reset) begin
      _T_2392_0 <= 1'h0;
    end else begin
      _T_2392_0 <= _T_2235;
    end
    if (reset) begin
      _T_2392_1 <= 1'h0;
    end else begin
      _T_2392_1 <= _T_2392_0;
    end
    if (reset) begin
      _T_2392_2 <= 1'h0;
    end else begin
      _T_2392_2 <= _T_2392_1;
    end
    if (reset) begin
      _T_2392_3 <= 1'h0;
    end else begin
      _T_2392_3 <= _T_2392_2;
    end
    if (reset) begin
      _T_2402_0 <= 1'h0;
    end else begin
      _T_2402_0 <= _T_2395;
    end
    if (reset) begin
      _T_2402_1 <= 1'h0;
    end else begin
      _T_2402_1 <= _T_2402_0;
    end
    if (reset) begin
      _T_2402_2 <= 1'h0;
    end else begin
      _T_2402_2 <= _T_2402_1;
    end
    if (reset) begin
      _T_2402_3 <= 1'h0;
    end else begin
      _T_2402_3 <= _T_2402_2;
    end
    if (reset) begin
      _T_2412_0 <= 1'h0;
    end else begin
      _T_2412_0 <= _T_155;
    end
    if (reset) begin
      _T_2412_1 <= 1'h0;
    end else begin
      _T_2412_1 <= _T_2412_0;
    end
    if (reset) begin
      _T_2412_2 <= 1'h0;
    end else begin
      _T_2412_2 <= _T_2412_1;
    end
    if (reset) begin
      _T_2412_3 <= 1'h0;
    end else begin
      _T_2412_3 <= _T_2412_2;
    end
    if (reset) begin
      _T_2422_0 <= 1'h0;
    end else begin
      _T_2422_0 <= _T_315;
    end
    if (reset) begin
      _T_2422_1 <= 1'h0;
    end else begin
      _T_2422_1 <= _T_2422_0;
    end
    if (reset) begin
      _T_2422_2 <= 1'h0;
    end else begin
      _T_2422_2 <= _T_2422_1;
    end
    if (reset) begin
      _T_2422_3 <= 1'h0;
    end else begin
      _T_2422_3 <= _T_2422_2;
    end
    if (reset) begin
      _T_2432_0 <= 1'h0;
    end else begin
      _T_2432_0 <= _T_475;
    end
    if (reset) begin
      _T_2432_1 <= 1'h0;
    end else begin
      _T_2432_1 <= _T_2432_0;
    end
    if (reset) begin
      _T_2432_2 <= 1'h0;
    end else begin
      _T_2432_2 <= _T_2432_1;
    end
    if (reset) begin
      _T_2432_3 <= 1'h0;
    end else begin
      _T_2432_3 <= _T_2432_2;
    end
    if (reset) begin
      _T_2442_0 <= 1'h0;
    end else begin
      _T_2442_0 <= _T_635;
    end
    if (reset) begin
      _T_2442_1 <= 1'h0;
    end else begin
      _T_2442_1 <= _T_2442_0;
    end
    if (reset) begin
      _T_2442_2 <= 1'h0;
    end else begin
      _T_2442_2 <= _T_2442_1;
    end
    if (reset) begin
      _T_2442_3 <= 1'h0;
    end else begin
      _T_2442_3 <= _T_2442_2;
    end
    if (reset) begin
      _T_2452_0 <= 1'h0;
    end else begin
      _T_2452_0 <= _T_795;
    end
    if (reset) begin
      _T_2452_1 <= 1'h0;
    end else begin
      _T_2452_1 <= _T_2452_0;
    end
    if (reset) begin
      _T_2452_2 <= 1'h0;
    end else begin
      _T_2452_2 <= _T_2452_1;
    end
    if (reset) begin
      _T_2452_3 <= 1'h0;
    end else begin
      _T_2452_3 <= _T_2452_2;
    end
    if (reset) begin
      _T_2462_0 <= 1'h0;
    end else begin
      _T_2462_0 <= _T_955;
    end
    if (reset) begin
      _T_2462_1 <= 1'h0;
    end else begin
      _T_2462_1 <= _T_2462_0;
    end
    if (reset) begin
      _T_2462_2 <= 1'h0;
    end else begin
      _T_2462_2 <= _T_2462_1;
    end
    if (reset) begin
      _T_2462_3 <= 1'h0;
    end else begin
      _T_2462_3 <= _T_2462_2;
    end
    if (reset) begin
      _T_2472_0 <= 1'h0;
    end else begin
      _T_2472_0 <= _T_1115;
    end
    if (reset) begin
      _T_2472_1 <= 1'h0;
    end else begin
      _T_2472_1 <= _T_2472_0;
    end
    if (reset) begin
      _T_2472_2 <= 1'h0;
    end else begin
      _T_2472_2 <= _T_2472_1;
    end
    if (reset) begin
      _T_2472_3 <= 1'h0;
    end else begin
      _T_2472_3 <= _T_2472_2;
    end
    if (reset) begin
      _T_2482_0 <= 1'h0;
    end else begin
      _T_2482_0 <= _T_1275;
    end
    if (reset) begin
      _T_2482_1 <= 1'h0;
    end else begin
      _T_2482_1 <= _T_2482_0;
    end
    if (reset) begin
      _T_2482_2 <= 1'h0;
    end else begin
      _T_2482_2 <= _T_2482_1;
    end
    if (reset) begin
      _T_2482_3 <= 1'h0;
    end else begin
      _T_2482_3 <= _T_2482_2;
    end
    if (reset) begin
      _T_2492_0 <= 1'h0;
    end else begin
      _T_2492_0 <= _T_1435;
    end
    if (reset) begin
      _T_2492_1 <= 1'h0;
    end else begin
      _T_2492_1 <= _T_2492_0;
    end
    if (reset) begin
      _T_2492_2 <= 1'h0;
    end else begin
      _T_2492_2 <= _T_2492_1;
    end
    if (reset) begin
      _T_2492_3 <= 1'h0;
    end else begin
      _T_2492_3 <= _T_2492_2;
    end
    if (reset) begin
      _T_2502_0 <= 1'h0;
    end else begin
      _T_2502_0 <= _T_1595;
    end
    if (reset) begin
      _T_2502_1 <= 1'h0;
    end else begin
      _T_2502_1 <= _T_2502_0;
    end
    if (reset) begin
      _T_2502_2 <= 1'h0;
    end else begin
      _T_2502_2 <= _T_2502_1;
    end
    if (reset) begin
      _T_2502_3 <= 1'h0;
    end else begin
      _T_2502_3 <= _T_2502_2;
    end
    if (reset) begin
      _T_2512_0 <= 1'h0;
    end else begin
      _T_2512_0 <= _T_1755;
    end
    if (reset) begin
      _T_2512_1 <= 1'h0;
    end else begin
      _T_2512_1 <= _T_2512_0;
    end
    if (reset) begin
      _T_2512_2 <= 1'h0;
    end else begin
      _T_2512_2 <= _T_2512_1;
    end
    if (reset) begin
      _T_2512_3 <= 1'h0;
    end else begin
      _T_2512_3 <= _T_2512_2;
    end
    if (reset) begin
      _T_2522_0 <= 1'h0;
    end else begin
      _T_2522_0 <= _T_1915;
    end
    if (reset) begin
      _T_2522_1 <= 1'h0;
    end else begin
      _T_2522_1 <= _T_2522_0;
    end
    if (reset) begin
      _T_2522_2 <= 1'h0;
    end else begin
      _T_2522_2 <= _T_2522_1;
    end
    if (reset) begin
      _T_2522_3 <= 1'h0;
    end else begin
      _T_2522_3 <= _T_2522_2;
    end
    if (reset) begin
      _T_2532_0 <= 1'h0;
    end else begin
      _T_2532_0 <= _T_2075;
    end
    if (reset) begin
      _T_2532_1 <= 1'h0;
    end else begin
      _T_2532_1 <= _T_2532_0;
    end
    if (reset) begin
      _T_2532_2 <= 1'h0;
    end else begin
      _T_2532_2 <= _T_2532_1;
    end
    if (reset) begin
      _T_2532_3 <= 1'h0;
    end else begin
      _T_2532_3 <= _T_2532_2;
    end
    if (reset) begin
      _T_2542_0 <= 1'h0;
    end else begin
      _T_2542_0 <= _T_2235;
    end
    if (reset) begin
      _T_2542_1 <= 1'h0;
    end else begin
      _T_2542_1 <= _T_2542_0;
    end
    if (reset) begin
      _T_2542_2 <= 1'h0;
    end else begin
      _T_2542_2 <= _T_2542_1;
    end
    if (reset) begin
      _T_2542_3 <= 1'h0;
    end else begin
      _T_2542_3 <= _T_2542_2;
    end
    if (reset) begin
      _T_2552_0 <= 1'h0;
    end else begin
      _T_2552_0 <= _T_2395;
    end
    if (reset) begin
      _T_2552_1 <= 1'h0;
    end else begin
      _T_2552_1 <= _T_2552_0;
    end
    if (reset) begin
      _T_2552_2 <= 1'h0;
    end else begin
      _T_2552_2 <= _T_2552_1;
    end
    if (reset) begin
      _T_2552_3 <= 1'h0;
    end else begin
      _T_2552_3 <= _T_2552_2;
    end
    if (reset) begin
      _T_2562_0 <= 1'h0;
    end else begin
      _T_2562_0 <= _T_2555;
    end
    if (reset) begin
      _T_2562_1 <= 1'h0;
    end else begin
      _T_2562_1 <= _T_2562_0;
    end
    if (reset) begin
      _T_2562_2 <= 1'h0;
    end else begin
      _T_2562_2 <= _T_2562_1;
    end
    if (reset) begin
      _T_2562_3 <= 1'h0;
    end else begin
      _T_2562_3 <= _T_2562_2;
    end
    if (reset) begin
      _T_2575_0 <= 1'h0;
    end else begin
      _T_2575_0 <= _T_2570;
    end
    if (reset) begin
      _T_2575_1 <= 1'h0;
    end else begin
      _T_2575_1 <= _T_2575_0;
    end
    if (reset) begin
      _T_2575_2 <= 1'h0;
    end else begin
      _T_2575_2 <= _T_2575_1;
    end
    if (reset) begin
      _T_2584_0 <= 1'h0;
    end else begin
      _T_2584_0 <= _T_2579;
    end
    if (reset) begin
      _T_2584_1 <= 1'h0;
    end else begin
      _T_2584_1 <= _T_2584_0;
    end
    if (reset) begin
      _T_2584_2 <= 1'h0;
    end else begin
      _T_2584_2 <= _T_2584_1;
    end
    if (reset) begin
      _T_2593_0 <= 1'h0;
    end else begin
      _T_2593_0 <= _T_2588;
    end
    if (reset) begin
      _T_2593_1 <= 1'h0;
    end else begin
      _T_2593_1 <= _T_2593_0;
    end
    if (reset) begin
      _T_2593_2 <= 1'h0;
    end else begin
      _T_2593_2 <= _T_2593_1;
    end
    if (reset) begin
      _T_2602_0 <= 1'h0;
    end else begin
      _T_2602_0 <= _T_2597;
    end
    if (reset) begin
      _T_2602_1 <= 1'h0;
    end else begin
      _T_2602_1 <= _T_2602_0;
    end
    if (reset) begin
      _T_2602_2 <= 1'h0;
    end else begin
      _T_2602_2 <= _T_2602_1;
    end
    if (reset) begin
      _T_2611_0 <= 1'h0;
    end else begin
      _T_2611_0 <= _T_2606;
    end
    if (reset) begin
      _T_2611_1 <= 1'h0;
    end else begin
      _T_2611_1 <= _T_2611_0;
    end
    if (reset) begin
      _T_2611_2 <= 1'h0;
    end else begin
      _T_2611_2 <= _T_2611_1;
    end
    if (reset) begin
      _T_2620_0 <= 1'h0;
    end else begin
      _T_2620_0 <= _T_2615;
    end
    if (reset) begin
      _T_2620_1 <= 1'h0;
    end else begin
      _T_2620_1 <= _T_2620_0;
    end
    if (reset) begin
      _T_2620_2 <= 1'h0;
    end else begin
      _T_2620_2 <= _T_2620_1;
    end
    if (reset) begin
      _T_2629_0 <= 1'h0;
    end else begin
      _T_2629_0 <= _T_2624;
    end
    if (reset) begin
      _T_2629_1 <= 1'h0;
    end else begin
      _T_2629_1 <= _T_2629_0;
    end
    if (reset) begin
      _T_2629_2 <= 1'h0;
    end else begin
      _T_2629_2 <= _T_2629_1;
    end
    if (reset) begin
      _T_2638_0 <= 1'h0;
    end else begin
      _T_2638_0 <= _T_2633;
    end
    if (reset) begin
      _T_2638_1 <= 1'h0;
    end else begin
      _T_2638_1 <= _T_2638_0;
    end
    if (reset) begin
      _T_2638_2 <= 1'h0;
    end else begin
      _T_2638_2 <= _T_2638_1;
    end
    if (reset) begin
      _T_2647_0 <= 1'h0;
    end else begin
      _T_2647_0 <= _T_2642;
    end
    if (reset) begin
      _T_2647_1 <= 1'h0;
    end else begin
      _T_2647_1 <= _T_2647_0;
    end
    if (reset) begin
      _T_2647_2 <= 1'h0;
    end else begin
      _T_2647_2 <= _T_2647_1;
    end
    if (reset) begin
      _T_2656_0 <= 1'h0;
    end else begin
      _T_2656_0 <= _T_2651;
    end
    if (reset) begin
      _T_2656_1 <= 1'h0;
    end else begin
      _T_2656_1 <= _T_2656_0;
    end
    if (reset) begin
      _T_2656_2 <= 1'h0;
    end else begin
      _T_2656_2 <= _T_2656_1;
    end
    if (reset) begin
      _T_2665_0 <= 1'h0;
    end else begin
      _T_2665_0 <= _T_2660;
    end
    if (reset) begin
      _T_2665_1 <= 1'h0;
    end else begin
      _T_2665_1 <= _T_2665_0;
    end
    if (reset) begin
      _T_2665_2 <= 1'h0;
    end else begin
      _T_2665_2 <= _T_2665_1;
    end
    if (reset) begin
      _T_2674_0 <= 1'h0;
    end else begin
      _T_2674_0 <= _T_2669;
    end
    if (reset) begin
      _T_2674_1 <= 1'h0;
    end else begin
      _T_2674_1 <= _T_2674_0;
    end
    if (reset) begin
      _T_2674_2 <= 1'h0;
    end else begin
      _T_2674_2 <= _T_2674_1;
    end
    if (reset) begin
      _T_2683_0 <= 1'h0;
    end else begin
      _T_2683_0 <= _T_2678;
    end
    if (reset) begin
      _T_2683_1 <= 1'h0;
    end else begin
      _T_2683_1 <= _T_2683_0;
    end
    if (reset) begin
      _T_2683_2 <= 1'h0;
    end else begin
      _T_2683_2 <= _T_2683_1;
    end
    if (reset) begin
      _T_2692_0 <= 1'h0;
    end else begin
      _T_2692_0 <= _T_2687;
    end
    if (reset) begin
      _T_2692_1 <= 1'h0;
    end else begin
      _T_2692_1 <= _T_2692_0;
    end
    if (reset) begin
      _T_2692_2 <= 1'h0;
    end else begin
      _T_2692_2 <= _T_2692_1;
    end
    if (reset) begin
      _T_2701_0 <= 1'h0;
    end else begin
      _T_2701_0 <= _T_2696;
    end
    if (reset) begin
      _T_2701_1 <= 1'h0;
    end else begin
      _T_2701_1 <= _T_2701_0;
    end
    if (reset) begin
      _T_2701_2 <= 1'h0;
    end else begin
      _T_2701_2 <= _T_2701_1;
    end
    if (reset) begin
      _T_2710_0 <= 1'h0;
    end else begin
      _T_2710_0 <= _T_2705;
    end
    if (reset) begin
      _T_2710_1 <= 1'h0;
    end else begin
      _T_2710_1 <= _T_2710_0;
    end
    if (reset) begin
      _T_2710_2 <= 1'h0;
    end else begin
      _T_2710_2 <= _T_2710_1;
    end
    if (reset) begin
      _T_2712_0 <= 1'h0;
    end else begin
      _T_2712_0 <= io_exec_valid;
    end
    if (reset) begin
      _T_2712_1 <= 1'h0;
    end else begin
      _T_2712_1 <= _T_2712_0;
    end
    if (reset) begin
      _T_2712_2 <= 1'h0;
    end else begin
      _T_2712_2 <= _T_2712_1;
    end
    if (reset) begin
      _T_2712_3 <= 1'h0;
    end else begin
      _T_2712_3 <= _T_2712_2;
    end
    if (reset) begin
      _T_2712_4 <= 1'h0;
    end else begin
      _T_2712_4 <= _T_2712_3;
    end
    if (reset) begin
      _T_2712_5 <= 1'h0;
    end else begin
      _T_2712_5 <= _T_2712_4;
    end
    if (reset) begin
      _T_2712_6 <= 1'h0;
    end else begin
      _T_2712_6 <= _T_2712_5;
    end
    if (reset) begin
      _T_2712_7 <= 1'h0;
    end else begin
      _T_2712_7 <= _T_2712_6;
    end
    if (reset) begin
      _T_2712_8 <= 1'h0;
    end else begin
      _T_2712_8 <= _T_2712_7;
    end
    if (reset) begin
      _T_2712_9 <= 1'h0;
    end else begin
      _T_2712_9 <= _T_2712_8;
    end
    if (reset) begin
      _T_2712_10 <= 1'h0;
    end else begin
      _T_2712_10 <= _T_2712_9;
    end
    if (reset) begin
      _T_2712_11 <= 1'h0;
    end else begin
      _T_2712_11 <= _T_2712_10;
    end
    if (reset) begin
      _T_2712_12 <= 1'h0;
    end else begin
      _T_2712_12 <= _T_2712_11;
    end
    if (reset) begin
      _T_2712_13 <= 1'h0;
    end else begin
      _T_2712_13 <= _T_2712_12;
    end
    if (reset) begin
      _T_2712_14 <= 1'h0;
    end else begin
      _T_2712_14 <= _T_2712_13;
    end
    if (reset) begin
      _T_2712_15 <= 1'h0;
    end else begin
      _T_2712_15 <= _T_2712_14;
    end
    if (reset) begin
      _T_2712_16 <= 1'h0;
    end else begin
      _T_2712_16 <= _T_2712_15;
    end
    if (reset) begin
      _T_2712_17 <= 1'h0;
    end else begin
      _T_2712_17 <= _T_2712_16;
    end
    if (reset) begin
      _T_2712_18 <= 1'h0;
    end else begin
      _T_2712_18 <= _T_2712_17;
    end
    if (reset) begin
      _T_2712_19 <= 1'h0;
    end else begin
      _T_2712_19 <= _T_2712_18;
    end
    if (reset) begin
      _T_2712_20 <= 1'h0;
    end else begin
      _T_2712_20 <= _T_2712_19;
    end
    if (reset) begin
      _T_2712_21 <= 1'h0;
    end else begin
      _T_2712_21 <= _T_2712_20;
    end
    if (reset) begin
      _T_2712_22 <= 1'h0;
    end else begin
      _T_2712_22 <= _T_2712_21;
    end
    if (reset) begin
      _T_2712_23 <= 1'h0;
    end else begin
      _T_2712_23 <= _T_2712_22;
    end
    if (reset) begin
      _T_2712_24 <= 1'h0;
    end else begin
      _T_2712_24 <= _T_2712_23;
    end
    if (reset) begin
      _T_2712_25 <= 1'h0;
    end else begin
      _T_2712_25 <= _T_2712_24;
    end
    if (reset) begin
      _T_2712_26 <= 1'h0;
    end else begin
      _T_2712_26 <= _T_2712_25;
    end
    if (reset) begin
      _T_2712_27 <= 1'h0;
    end else begin
      _T_2712_27 <= _T_2712_26;
    end
    if (reset) begin
      _T_2712_28 <= 1'h0;
    end else begin
      _T_2712_28 <= _T_2712_27;
    end
    if (reset) begin
      _T_2712_29 <= 1'h0;
    end else begin
      _T_2712_29 <= _T_2712_28;
    end
    if (reset) begin
      _T_2712_30 <= 1'h0;
    end else begin
      _T_2712_30 <= _T_2712_29;
    end
    if (reset) begin
      _T_2712_31 <= 1'h0;
    end else begin
      _T_2712_31 <= _T_2712_30;
    end
    if (reset) begin
      _T_2712_32 <= 1'h0;
    end else begin
      _T_2712_32 <= _T_2712_31;
    end
    if (reset) begin
      _T_2712_33 <= 1'h0;
    end else begin
      _T_2712_33 <= _T_2712_32;
    end
    if (reset) begin
      _T_2712_34 <= 1'h0;
    end else begin
      _T_2712_34 <= _T_2712_33;
    end
    if (reset) begin
      _T_2712_35 <= 1'h0;
    end else begin
      _T_2712_35 <= _T_2712_34;
    end
    if (reset) begin
      _T_2712_36 <= 1'h0;
    end else begin
      _T_2712_36 <= _T_2712_35;
    end
    if (reset) begin
      _T_2712_37 <= 1'h0;
    end else begin
      _T_2712_37 <= _T_2712_36;
    end
    if (reset) begin
      _T_2712_38 <= 1'h0;
    end else begin
      _T_2712_38 <= _T_2712_37;
    end
    if (reset) begin
      _T_2712_39 <= 1'h0;
    end else begin
      _T_2712_39 <= _T_2712_38;
    end
    if (reset) begin
      _T_2712_40 <= 1'h0;
    end else begin
      _T_2712_40 <= _T_2712_39;
    end
    if (reset) begin
      _T_2712_41 <= 1'h0;
    end else begin
      _T_2712_41 <= _T_2712_40;
    end
    if (reset) begin
      _T_2712_42 <= 1'h0;
    end else begin
      _T_2712_42 <= _T_2712_41;
    end
    if (reset) begin
      _T_2712_43 <= 1'h0;
    end else begin
      _T_2712_43 <= _T_2712_42;
    end
    if (reset) begin
      _T_2712_44 <= 1'h0;
    end else begin
      _T_2712_44 <= _T_2712_43;
    end
    if (reset) begin
      _T_2712_45 <= 1'h0;
    end else begin
      _T_2712_45 <= _T_2712_44;
    end
    if (reset) begin
      _T_2712_46 <= 1'h0;
    end else begin
      _T_2712_46 <= _T_2712_45;
    end
    if (reset) begin
      _T_2712_47 <= 1'h0;
    end else begin
      _T_2712_47 <= _T_2712_46;
    end
    if (reset) begin
      _T_2712_48 <= 1'h0;
    end else begin
      _T_2712_48 <= _T_2712_47;
    end
    if (reset) begin
      _T_2712_49 <= 1'h0;
    end else begin
      _T_2712_49 <= _T_2712_48;
    end
    if (reset) begin
      _T_2712_50 <= 1'h0;
    end else begin
      _T_2712_50 <= _T_2712_49;
    end
    if (reset) begin
      _T_2712_51 <= 1'h0;
    end else begin
      _T_2712_51 <= _T_2712_50;
    end
    if (reset) begin
      _T_2712_52 <= 1'h0;
    end else begin
      _T_2712_52 <= _T_2712_51;
    end
    if (reset) begin
      _T_2712_53 <= 1'h0;
    end else begin
      _T_2712_53 <= _T_2712_52;
    end
    if (reset) begin
      _T_2712_54 <= 1'h0;
    end else begin
      _T_2712_54 <= _T_2712_53;
    end
    if (reset) begin
      _T_2712_55 <= 1'h0;
    end else begin
      _T_2712_55 <= _T_2712_54;
    end
    if (reset) begin
      _T_2712_56 <= 1'h0;
    end else begin
      _T_2712_56 <= _T_2712_55;
    end
    if (reset) begin
      _T_2712_57 <= 1'h0;
    end else begin
      _T_2712_57 <= _T_2712_56;
    end
    if (reset) begin
      _T_2712_58 <= 1'h0;
    end else begin
      _T_2712_58 <= _T_2712_57;
    end
    if (reset) begin
      _T_2712_59 <= 1'h0;
    end else begin
      _T_2712_59 <= _T_2712_58;
    end
    if (reset) begin
      _T_2712_60 <= 1'h0;
    end else begin
      _T_2712_60 <= _T_2712_59;
    end
    if (reset) begin
      _T_2712_61 <= 1'h0;
    end else begin
      _T_2712_61 <= _T_2712_60;
    end
    if (reset) begin
      _T_2712_62 <= 1'h0;
    end else begin
      _T_2712_62 <= _T_2712_61;
    end
    if (reset) begin
      _T_2712_63 <= 1'h0;
    end else begin
      _T_2712_63 <= _T_2712_62;
    end
    if (reset) begin
      _T_2712_64 <= 1'h0;
    end else begin
      _T_2712_64 <= _T_2712_63;
    end
    if (reset) begin
      _T_2712_65 <= 1'h0;
    end else begin
      _T_2712_65 <= _T_2712_64;
    end
    if (reset) begin
      _T_2712_66 <= 1'h0;
    end else begin
      _T_2712_66 <= _T_2712_65;
    end
    if (reset) begin
      _T_2712_67 <= 1'h0;
    end else begin
      _T_2712_67 <= _T_2712_66;
    end
    if (reset) begin
      _T_2712_68 <= 1'h0;
    end else begin
      _T_2712_68 <= _T_2712_67;
    end
    if (reset) begin
      _T_2712_69 <= 1'h0;
    end else begin
      _T_2712_69 <= _T_2712_68;
    end
    if (reset) begin
      _T_2712_70 <= 1'h0;
    end else begin
      _T_2712_70 <= _T_2712_69;
    end
    if (reset) begin
      _T_2712_71 <= 1'h0;
    end else begin
      _T_2712_71 <= _T_2712_70;
    end
    if (reset) begin
      _T_2712_72 <= 1'h0;
    end else begin
      _T_2712_72 <= _T_2712_71;
    end
    if (reset) begin
      _T_2712_73 <= 1'h0;
    end else begin
      _T_2712_73 <= _T_2712_72;
    end
    if (reset) begin
      _T_2712_74 <= 1'h0;
    end else begin
      _T_2712_74 <= _T_2712_73;
    end
    if (reset) begin
      _T_2712_75 <= 1'h0;
    end else begin
      _T_2712_75 <= _T_2712_74;
    end
    if (reset) begin
      _T_2712_76 <= 1'h0;
    end else begin
      _T_2712_76 <= _T_2712_75;
    end
    if (reset) begin
      _T_2712_77 <= 1'h0;
    end else begin
      _T_2712_77 <= _T_2712_76;
    end
    if (reset) begin
      _T_2712_78 <= 1'h0;
    end else begin
      _T_2712_78 <= _T_2712_77;
    end
    if (reset) begin
      _T_2712_79 <= 1'h0;
    end else begin
      _T_2712_79 <= _T_2712_78;
    end
    if (reset) begin
      _T_2712_80 <= 1'h0;
    end else begin
      _T_2712_80 <= _T_2712_79;
    end
    if (reset) begin
      _T_2712_81 <= 1'h0;
    end else begin
      _T_2712_81 <= _T_2712_80;
    end
    if (reset) begin
      _T_2712_82 <= 1'h0;
    end else begin
      _T_2712_82 <= _T_2712_81;
    end
    if (reset) begin
      _T_2712_83 <= 1'h0;
    end else begin
      _T_2712_83 <= _T_2712_82;
    end
    if (reset) begin
      _T_2712_84 <= 1'h0;
    end else begin
      _T_2712_84 <= _T_2712_83;
    end
    if (reset) begin
      _T_2712_85 <= 1'h0;
    end else begin
      _T_2712_85 <= _T_2712_84;
    end
    if (reset) begin
      _T_2712_86 <= 1'h0;
    end else begin
      _T_2712_86 <= _T_2712_85;
    end
    if (reset) begin
      _T_2712_87 <= 1'h0;
    end else begin
      _T_2712_87 <= _T_2712_86;
    end
    if (reset) begin
      _T_2712_88 <= 1'h0;
    end else begin
      _T_2712_88 <= _T_2712_87;
    end
    if (reset) begin
      _T_2712_89 <= 1'h0;
    end else begin
      _T_2712_89 <= _T_2712_88;
    end
    if (reset) begin
      _T_2712_90 <= 1'h0;
    end else begin
      _T_2712_90 <= _T_2712_89;
    end
    if (reset) begin
      _T_2712_91 <= 1'h0;
    end else begin
      _T_2712_91 <= _T_2712_90;
    end
    if (reset) begin
      _T_2712_92 <= 1'h0;
    end else begin
      _T_2712_92 <= _T_2712_91;
    end
    if (reset) begin
      _T_2712_93 <= 1'h0;
    end else begin
      _T_2712_93 <= _T_2712_92;
    end
    if (reset) begin
      _T_2712_94 <= 1'h0;
    end else begin
      _T_2712_94 <= _T_2712_93;
    end
    if (reset) begin
      _T_2712_95 <= 1'h0;
    end else begin
      _T_2712_95 <= _T_2712_94;
    end
    if (reset) begin
      _T_2712_96 <= 1'h0;
    end else begin
      _T_2712_96 <= _T_2712_95;
    end
    if (reset) begin
      _T_2712_97 <= 1'h0;
    end else begin
      _T_2712_97 <= _T_2712_96;
    end
    if (reset) begin
      _T_2712_98 <= 1'h0;
    end else begin
      _T_2712_98 <= _T_2712_97;
    end
    if (reset) begin
      _T_2712_99 <= 1'h0;
    end else begin
      _T_2712_99 <= _T_2712_98;
    end
    if (reset) begin
      _T_2712_100 <= 1'h0;
    end else begin
      _T_2712_100 <= _T_2712_99;
    end
    if (reset) begin
      _T_2712_101 <= 1'h0;
    end else begin
      _T_2712_101 <= _T_2712_100;
    end
    if (reset) begin
      _T_2712_102 <= 1'h0;
    end else begin
      _T_2712_102 <= _T_2712_101;
    end
    if (reset) begin
      _T_2712_103 <= 1'h0;
    end else begin
      _T_2712_103 <= _T_2712_102;
    end
    if (reset) begin
      _T_2712_104 <= 1'h0;
    end else begin
      _T_2712_104 <= _T_2712_103;
    end
    if (reset) begin
      _T_2712_105 <= 1'h0;
    end else begin
      _T_2712_105 <= _T_2712_104;
    end
    if (reset) begin
      _T_2712_106 <= 1'h0;
    end else begin
      _T_2712_106 <= _T_2712_105;
    end
    if (reset) begin
      _T_2712_107 <= 1'h0;
    end else begin
      _T_2712_107 <= _T_2712_106;
    end
    if (reset) begin
      _T_2712_108 <= 1'h0;
    end else begin
      _T_2712_108 <= _T_2712_107;
    end
    if (reset) begin
      _T_2712_109 <= 1'h0;
    end else begin
      _T_2712_109 <= _T_2712_108;
    end
    if (reset) begin
      _T_2712_110 <= 1'h0;
    end else begin
      _T_2712_110 <= _T_2712_109;
    end
    if (reset) begin
      _T_2712_111 <= 1'h0;
    end else begin
      _T_2712_111 <= _T_2712_110;
    end
    if (reset) begin
      _T_2712_112 <= 1'h0;
    end else begin
      _T_2712_112 <= _T_2712_111;
    end
    if (reset) begin
      _T_2712_113 <= 1'h0;
    end else begin
      _T_2712_113 <= _T_2712_112;
    end
    if (reset) begin
      _T_2712_114 <= 1'h0;
    end else begin
      _T_2712_114 <= _T_2712_113;
    end
    if (reset) begin
      _T_2712_115 <= 1'h0;
    end else begin
      _T_2712_115 <= _T_2712_114;
    end
    if (reset) begin
      _T_2712_116 <= 1'h0;
    end else begin
      _T_2712_116 <= _T_2712_115;
    end
    if (reset) begin
      _T_2712_117 <= 1'h0;
    end else begin
      _T_2712_117 <= _T_2712_116;
    end
    if (reset) begin
      _T_2712_118 <= 1'h0;
    end else begin
      _T_2712_118 <= _T_2712_117;
    end
    if (reset) begin
      _T_2712_119 <= 1'h0;
    end else begin
      _T_2712_119 <= _T_2712_118;
    end
    if (reset) begin
      _T_2712_120 <= 1'h0;
    end else begin
      _T_2712_120 <= _T_2712_119;
    end
    if (reset) begin
      _T_2712_121 <= 1'h0;
    end else begin
      _T_2712_121 <= _T_2712_120;
    end
    if (reset) begin
      _T_2712_122 <= 1'h0;
    end else begin
      _T_2712_122 <= _T_2712_121;
    end
    if (reset) begin
      _T_2712_123 <= 1'h0;
    end else begin
      _T_2712_123 <= _T_2712_122;
    end
    if (reset) begin
      _T_2712_124 <= 1'h0;
    end else begin
      _T_2712_124 <= _T_2712_123;
    end
    if (reset) begin
      _T_2712_125 <= 1'h0;
    end else begin
      _T_2712_125 <= _T_2712_124;
    end
    if (reset) begin
      _T_2712_126 <= 1'h0;
    end else begin
      _T_2712_126 <= _T_2712_125;
    end
    if (reset) begin
      _T_2712_127 <= 1'h0;
    end else begin
      _T_2712_127 <= _T_2712_126;
    end
    if (reset) begin
      _T_2712_128 <= 1'h0;
    end else begin
      _T_2712_128 <= _T_2712_127;
    end
    if (reset) begin
      _T_2712_129 <= 1'h0;
    end else begin
      _T_2712_129 <= _T_2712_128;
    end
    if (reset) begin
      _T_2712_130 <= 1'h0;
    end else begin
      _T_2712_130 <= _T_2712_129;
    end
    if (reset) begin
      _T_2712_131 <= 1'h0;
    end else begin
      _T_2712_131 <= _T_2712_130;
    end
    if (reset) begin
      _T_2712_132 <= 1'h0;
    end else begin
      _T_2712_132 <= _T_2712_131;
    end
    if (reset) begin
      _T_2712_133 <= 1'h0;
    end else begin
      _T_2712_133 <= _T_2712_132;
    end
    if (reset) begin
      _T_2712_134 <= 1'h0;
    end else begin
      _T_2712_134 <= _T_2712_133;
    end
    if (reset) begin
      _T_2712_135 <= 1'h0;
    end else begin
      _T_2712_135 <= _T_2712_134;
    end
    if (reset) begin
      _T_2712_136 <= 1'h0;
    end else begin
      _T_2712_136 <= _T_2712_135;
    end
    if (reset) begin
      _T_2712_137 <= 1'h0;
    end else begin
      _T_2712_137 <= _T_2712_136;
    end
    if (reset) begin
      _T_2712_138 <= 1'h0;
    end else begin
      _T_2712_138 <= _T_2712_137;
    end
    if (reset) begin
      _T_2712_139 <= 1'h0;
    end else begin
      _T_2712_139 <= _T_2712_138;
    end
    if (reset) begin
      _T_2712_140 <= 1'h0;
    end else begin
      _T_2712_140 <= _T_2712_139;
    end
    if (reset) begin
      _T_2712_141 <= 1'h0;
    end else begin
      _T_2712_141 <= _T_2712_140;
    end
    if (reset) begin
      _T_2712_142 <= 1'h0;
    end else begin
      _T_2712_142 <= _T_2712_141;
    end
    if (reset) begin
      _T_2712_143 <= 1'h0;
    end else begin
      _T_2712_143 <= _T_2712_142;
    end
    if (reset) begin
      _T_2712_144 <= 1'h0;
    end else begin
      _T_2712_144 <= _T_2712_143;
    end
    if (reset) begin
      _T_2712_145 <= 1'h0;
    end else begin
      _T_2712_145 <= _T_2712_144;
    end
    if (reset) begin
      _T_2712_146 <= 1'h0;
    end else begin
      _T_2712_146 <= _T_2712_145;
    end
    if (reset) begin
      _T_2712_147 <= 1'h0;
    end else begin
      _T_2712_147 <= _T_2712_146;
    end
    if (reset) begin
      _T_2712_148 <= 1'h0;
    end else begin
      _T_2712_148 <= _T_2712_147;
    end
    if (reset) begin
      _T_2712_149 <= 1'h0;
    end else begin
      _T_2712_149 <= _T_2712_148;
    end
    if (reset) begin
      _T_2712_150 <= 1'h0;
    end else begin
      _T_2712_150 <= _T_2712_149;
    end
    if (reset) begin
      _T_2712_151 <= 1'h0;
    end else begin
      _T_2712_151 <= _T_2712_150;
    end
    if (reset) begin
      _T_2712_152 <= 1'h0;
    end else begin
      _T_2712_152 <= _T_2712_151;
    end
    if (reset) begin
      _T_2712_153 <= 1'h0;
    end else begin
      _T_2712_153 <= _T_2712_152;
    end
    if (reset) begin
      _T_2712_154 <= 1'h0;
    end else begin
      _T_2712_154 <= _T_2712_153;
    end
    if (reset) begin
      _T_2712_155 <= 1'h0;
    end else begin
      _T_2712_155 <= _T_2712_154;
    end
    if (reset) begin
      _T_2712_156 <= 1'h0;
    end else begin
      _T_2712_156 <= _T_2712_155;
    end
    if (reset) begin
      _T_2712_157 <= 1'h0;
    end else begin
      _T_2712_157 <= _T_2712_156;
    end
    if (reset) begin
      _T_2712_158 <= 1'h0;
    end else begin
      _T_2712_158 <= _T_2712_157;
    end
    if (reset) begin
      _T_2712_159 <= 1'h0;
    end else begin
      _T_2712_159 <= _T_2712_158;
    end
    if (reset) begin
      _T_2712_160 <= 1'h0;
    end else begin
      _T_2712_160 <= _T_2712_159;
    end
    if (reset) begin
      _T_2712_161 <= 1'h0;
    end else begin
      _T_2712_161 <= _T_2712_160;
    end
    if (reset) begin
      _T_2712_162 <= 1'h0;
    end else begin
      _T_2712_162 <= _T_2712_161;
    end
    if (reset) begin
      _T_2712_163 <= 1'h0;
    end else begin
      _T_2712_163 <= _T_2712_162;
    end
    if (reset) begin
      _T_2712_164 <= 1'h0;
    end else begin
      _T_2712_164 <= _T_2712_163;
    end
    if (reset) begin
      _T_2712_165 <= 1'h0;
    end else begin
      _T_2712_165 <= _T_2712_164;
    end
    if (reset) begin
      _T_2712_166 <= 1'h0;
    end else begin
      _T_2712_166 <= _T_2712_165;
    end
    if (reset) begin
      _T_2712_167 <= 1'h0;
    end else begin
      _T_2712_167 <= _T_2712_166;
    end
    if (reset) begin
      _T_2712_168 <= 1'h0;
    end else begin
      _T_2712_168 <= _T_2712_167;
    end
    if (reset) begin
      _T_2712_169 <= 1'h0;
    end else begin
      _T_2712_169 <= _T_2712_168;
    end
    if (reset) begin
      _T_2712_170 <= 1'h0;
    end else begin
      _T_2712_170 <= _T_2712_169;
    end
    if (reset) begin
      _T_2712_171 <= 1'h0;
    end else begin
      _T_2712_171 <= _T_2712_170;
    end
    if (reset) begin
      _T_2712_172 <= 1'h0;
    end else begin
      _T_2712_172 <= _T_2712_171;
    end
    if (reset) begin
      _T_2712_173 <= 1'h0;
    end else begin
      _T_2712_173 <= _T_2712_172;
    end
    if (reset) begin
      _T_2712_174 <= 1'h0;
    end else begin
      _T_2712_174 <= _T_2712_173;
    end
    if (reset) begin
      _T_2712_175 <= 1'h0;
    end else begin
      _T_2712_175 <= _T_2712_174;
    end
    if (reset) begin
      _T_2712_176 <= 1'h0;
    end else begin
      _T_2712_176 <= _T_2712_175;
    end
    if (reset) begin
      _T_2712_177 <= 1'h0;
    end else begin
      _T_2712_177 <= _T_2712_176;
    end
    if (reset) begin
      _T_2712_178 <= 1'h0;
    end else begin
      _T_2712_178 <= _T_2712_177;
    end
    if (reset) begin
      _T_2712_179 <= 1'h0;
    end else begin
      _T_2712_179 <= _T_2712_178;
    end
  end
endmodule
